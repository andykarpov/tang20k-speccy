--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.11 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Mon Jun 19 23:35:58 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(15 downto 0)
    );
end Gowin_pROM;

architecture Behavioral of Gowin_pROM is

    signal lut_f_0: std_logic;
    signal lut_f_1: std_logic;
    signal lut_f_2: std_logic;
    signal lut_f_3: std_logic;
    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_dout: std_logic_vector(0 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout: std_logic_vector(0 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout: std_logic_vector(0 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout: std_logic_vector(0 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout: std_logic_vector(1 downto 1);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout: std_logic_vector(1 downto 1);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout: std_logic_vector(1 downto 1);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout: std_logic_vector(1 downto 1);
    signal prom_inst_8_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_8_dout: std_logic_vector(2 downto 2);
    signal prom_inst_9_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_9_dout: std_logic_vector(2 downto 2);
    signal prom_inst_10_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_10_dout: std_logic_vector(2 downto 2);
    signal prom_inst_11_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_11_dout: std_logic_vector(2 downto 2);
    signal prom_inst_12_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_12_dout: std_logic_vector(3 downto 3);
    signal prom_inst_13_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_13_dout: std_logic_vector(3 downto 3);
    signal prom_inst_14_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_14_dout: std_logic_vector(3 downto 3);
    signal prom_inst_15_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_15_dout: std_logic_vector(3 downto 3);
    signal prom_inst_16_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_16_dout: std_logic_vector(4 downto 4);
    signal prom_inst_17_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_17_dout: std_logic_vector(4 downto 4);
    signal prom_inst_18_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_18_dout: std_logic_vector(4 downto 4);
    signal prom_inst_19_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_19_dout: std_logic_vector(4 downto 4);
    signal prom_inst_20_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_20_dout: std_logic_vector(5 downto 5);
    signal prom_inst_21_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_21_dout: std_logic_vector(5 downto 5);
    signal prom_inst_22_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_22_dout: std_logic_vector(5 downto 5);
    signal prom_inst_23_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_23_dout: std_logic_vector(5 downto 5);
    signal prom_inst_24_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_24_dout: std_logic_vector(6 downto 6);
    signal prom_inst_25_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_25_dout: std_logic_vector(6 downto 6);
    signal prom_inst_26_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_26_dout: std_logic_vector(6 downto 6);
    signal prom_inst_27_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_27_dout: std_logic_vector(6 downto 6);
    signal prom_inst_28_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_28_dout: std_logic_vector(7 downto 7);
    signal prom_inst_29_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_29_dout: std_logic_vector(7 downto 7);
    signal prom_inst_30_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_30_dout: std_logic_vector(7 downto 7);
    signal prom_inst_31_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_31_dout: std_logic_vector(7 downto 7);
    signal dff_q_0: std_logic;
    signal dff_q_1: std_logic;
    signal mux_o_0: std_logic;
    signal mux_o_1: std_logic;
    signal mux_o_3: std_logic;
    signal mux_o_4: std_logic;
    signal mux_o_6: std_logic;
    signal mux_o_7: std_logic;
    signal mux_o_9: std_logic;
    signal mux_o_10: std_logic;
    signal mux_o_12: std_logic;
    signal mux_o_13: std_logic;
    signal mux_o_15: std_logic;
    signal mux_o_16: std_logic;
    signal mux_o_18: std_logic;
    signal mux_o_19: std_logic;
    signal mux_o_21: std_logic;
    signal mux_o_22: std_logic;
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_8_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_9_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_10_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_11_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_12_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_13_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_14_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_15_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_16_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_17_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_18_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_19_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_20_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_21_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_22_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_23_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_24_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_25_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_26_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_27_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_28_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_29_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_30_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_31_DO_o: std_logic_vector(31 downto 0);

    -- component declaration
    component LUT3
        generic (
            INIT: in bit_vector := X"00"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic
        );
    end component;

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

    -- component declaration
    component DFFE
        port (
            Q: out std_logic;
            D: in std_logic;
            CLK: in std_logic;
            CE: in std_logic
        );
    end component;

    -- component declaration
    component MUX2
        port (
            O: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            S0: in std_logic
        );
    end component;

begin
    prom_inst_0_dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    prom_inst_1_dout(0) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    prom_inst_2_dout(0) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    prom_inst_3_dout(0) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    prom_inst_4_dout(1) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    prom_inst_5_dout(1) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    prom_inst_6_dout(1) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    prom_inst_7_dout(1) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;
    prom_inst_8_dout(2) <= prom_inst_8_DO_o(0);
    prom_inst_8_dout_w(30 downto 0) <= prom_inst_8_DO_o(31 downto 1) ;
    prom_inst_9_dout(2) <= prom_inst_9_DO_o(0);
    prom_inst_9_dout_w(30 downto 0) <= prom_inst_9_DO_o(31 downto 1) ;
    prom_inst_10_dout(2) <= prom_inst_10_DO_o(0);
    prom_inst_10_dout_w(30 downto 0) <= prom_inst_10_DO_o(31 downto 1) ;
    prom_inst_11_dout(2) <= prom_inst_11_DO_o(0);
    prom_inst_11_dout_w(30 downto 0) <= prom_inst_11_DO_o(31 downto 1) ;
    prom_inst_12_dout(3) <= prom_inst_12_DO_o(0);
    prom_inst_12_dout_w(30 downto 0) <= prom_inst_12_DO_o(31 downto 1) ;
    prom_inst_13_dout(3) <= prom_inst_13_DO_o(0);
    prom_inst_13_dout_w(30 downto 0) <= prom_inst_13_DO_o(31 downto 1) ;
    prom_inst_14_dout(3) <= prom_inst_14_DO_o(0);
    prom_inst_14_dout_w(30 downto 0) <= prom_inst_14_DO_o(31 downto 1) ;
    prom_inst_15_dout(3) <= prom_inst_15_DO_o(0);
    prom_inst_15_dout_w(30 downto 0) <= prom_inst_15_DO_o(31 downto 1) ;
    prom_inst_16_dout(4) <= prom_inst_16_DO_o(0);
    prom_inst_16_dout_w(30 downto 0) <= prom_inst_16_DO_o(31 downto 1) ;
    prom_inst_17_dout(4) <= prom_inst_17_DO_o(0);
    prom_inst_17_dout_w(30 downto 0) <= prom_inst_17_DO_o(31 downto 1) ;
    prom_inst_18_dout(4) <= prom_inst_18_DO_o(0);
    prom_inst_18_dout_w(30 downto 0) <= prom_inst_18_DO_o(31 downto 1) ;
    prom_inst_19_dout(4) <= prom_inst_19_DO_o(0);
    prom_inst_19_dout_w(30 downto 0) <= prom_inst_19_DO_o(31 downto 1) ;
    prom_inst_20_dout(5) <= prom_inst_20_DO_o(0);
    prom_inst_20_dout_w(30 downto 0) <= prom_inst_20_DO_o(31 downto 1) ;
    prom_inst_21_dout(5) <= prom_inst_21_DO_o(0);
    prom_inst_21_dout_w(30 downto 0) <= prom_inst_21_DO_o(31 downto 1) ;
    prom_inst_22_dout(5) <= prom_inst_22_DO_o(0);
    prom_inst_22_dout_w(30 downto 0) <= prom_inst_22_DO_o(31 downto 1) ;
    prom_inst_23_dout(5) <= prom_inst_23_DO_o(0);
    prom_inst_23_dout_w(30 downto 0) <= prom_inst_23_DO_o(31 downto 1) ;
    prom_inst_24_dout(6) <= prom_inst_24_DO_o(0);
    prom_inst_24_dout_w(30 downto 0) <= prom_inst_24_DO_o(31 downto 1) ;
    prom_inst_25_dout(6) <= prom_inst_25_DO_o(0);
    prom_inst_25_dout_w(30 downto 0) <= prom_inst_25_DO_o(31 downto 1) ;
    prom_inst_26_dout(6) <= prom_inst_26_DO_o(0);
    prom_inst_26_dout_w(30 downto 0) <= prom_inst_26_DO_o(31 downto 1) ;
    prom_inst_27_dout(6) <= prom_inst_27_DO_o(0);
    prom_inst_27_dout_w(30 downto 0) <= prom_inst_27_DO_o(31 downto 1) ;
    prom_inst_28_dout(7) <= prom_inst_28_DO_o(0);
    prom_inst_28_dout_w(30 downto 0) <= prom_inst_28_DO_o(31 downto 1) ;
    prom_inst_29_dout(7) <= prom_inst_29_DO_o(0);
    prom_inst_29_dout_w(30 downto 0) <= prom_inst_29_DO_o(31 downto 1) ;
    prom_inst_30_dout(7) <= prom_inst_30_DO_o(0);
    prom_inst_30_dout_w(30 downto 0) <= prom_inst_30_DO_o(31 downto 1) ;
    prom_inst_31_dout(7) <= prom_inst_31_DO_o(0);
    prom_inst_31_dout_w(30 downto 0) <= prom_inst_31_DO_o(31 downto 1) ;
    lut_inst_0 : LUT3
        generic map (
            INIT => X"02"
        )
        port map (
            F => lut_f_0,
            I0 => ce,
            I1 => ad(14),
            I2 => ad(15)
        );

    lut_inst_1 : LUT3
        generic map (
            INIT => X"08"
        )
        port map (
            F => lut_f_1,
            I0 => ce,
            I1 => ad(14),
            I2 => ad(15)
        );

    lut_inst_2 : LUT3
        generic map (
            INIT => X"20"
        )
        port map (
            F => lut_f_2,
            I0 => ce,
            I1 => ad(14),
            I2 => ad(15)
        );

    lut_inst_3 : LUT3
        generic map (
            INIT => X"80"
        )
        port map (
            F => lut_f_3,
            I0 => ce,
            I1 => ad(14),
            I2 => ad(15)
        );

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"352B1CB3ED3A7F8C2FFD607FCEBA3F08C9D6746F5995FADCAED4F9925B3995F3",
            INIT_RAM_01 => X"C99B2C66750F20C70263BBD92582182A4D582F00616B7CFB38D96C58229BA0F3",
            INIT_RAM_02 => X"9FE7EF999F9A613E9F3B221ADCF6DDED98B76C0411359EB7EA8B6CF7FD74DB39",
            INIT_RAM_03 => X"7FCC43F9E07FF5F7B7FFB7F43FFBAB30227FBFFADFCC229BB766E1E9BB1DD337",
            INIT_RAM_04 => X"F753B7D69DE33F40062F7CC2200006AB54007F9EFDFBFF36BBBB7D3F279EBD37",
            INIT_RAM_05 => X"53C5E2F714311FB17545D584A389DA684BD6EEC7C9727E7B3383FC3D9EA7FEEF",
            INIT_RAM_06 => X"9ABA0C567FB4EB3DDEEA2A35AA63453EE1ECF5A7F61F97F66CFD87E5F67B3F3E",
            INIT_RAM_07 => X"D17C7A32961E7478DFC018140683F37BFBFE7B72F66F6EFE9C173B3FFEF7ED26",
            INIT_RAM_08 => X"7AF88E7C0CFBEFB882E95651804688924D3403F93FED6BEF65D01BA62041FFF1",
            INIT_RAM_09 => X"C9178E5C66D2F7FFFFFCFEE7E9FBFFFFC0000002BFFFE3423CD538DC37AF239B",
            INIT_RAM_0A => X"41FD2ECFE6CD1FDBD37CEAE4EFCF5FD29B632B8FEFDE5C134AAADBB93D7CCE2C",
            INIT_RAM_0B => X"869FDDFB26DD2412BF6E5F332F3A3CF9FB9DA5E93C9FFEF6790F9E4EBFEFF7FC",
            INIT_RAM_0C => X"A3798FDB7FEB7A2ADA4B32ECFFE6AA889246099F76419D7208D39D7713DDA699",
            INIT_RAM_0D => X"526CB3DE4D9E4C9CB7F043828BC9F0AFDF2B7D5579BC7955454481DFF96EF8F0",
            INIT_RAM_0E => X"567B11080E43A75DC2158002801726EF841D647A75EF4449DD9B4696BE56749B",
            INIT_RAM_0F => X"DE014005764D523AEB374EA6D9B93FBAEB7A577E79C550E12F77762F3BF3DE09",
            INIT_RAM_10 => X"7757C5EF5492545AF576FEF75D9547FB1CD1CC50466056E8FE21E4FFF957CAC2",
            INIT_RAM_11 => X"5ADAD9E7CD3679F34D9A6CD379FBF26FCFD34EBAF4D3AEBFB2B2F795D5F5DFAB",
            INIT_RAM_12 => X"C357AC5224E91FBDDDAE6B91DCECD2668B1AFDFFFEEF7F4F7771524947BF65B2",
            INIT_RAM_13 => X"D0CBD11A22D0918161E9EFBA475FEEF342EFF7DDEFE7DFE9458C4FBF5BBE2E42",
            INIT_RAM_14 => X"DF7FAC98E34D5BAA0CD72E07DC6327FFDED8038DFFD8C9FFCC42E02BBE5EBE58",
            INIT_RAM_15 => X"89A70D55A17318A78ADD8BEF925534BC63257FB0D93EBF26FFAFAFD64F58CEDB",
            INIT_RAM_16 => X"674DD6BF7772BBFB7271F17BF7E9F0D04A728DC32DBD3A51CB83C8CECC468AEE",
            INIT_RAM_17 => X"EBF4D5555687F564A6BD5AE5FF3CB3F1E7F8EB559FCAA93B5236356090155131",
            INIT_RAM_18 => X"4132D95333C70B6F7E97BAD1336E66964FF55131FA52BB34E7D3FF91738E9DA8",
            INIT_RAM_19 => X"CF9A6CF3FD3FC6569BA7CFDECF3D1ACED3C7A3C7FBE7F6F3DDE1A9CF8DBADA3D",
            INIT_RAM_1A => X"F9E1EBDFC9FE79D006BEFC5EDE3FFF82FB4B22FA4DE351F4D3AEB9A6CF3E69B3",
            INIT_RAM_1B => X"AE555BD5B0D2D717BD367B0D9EEAB6ACF9FD1E95AC97F23B31BFF2774B31BA1F",
            INIT_RAM_1C => X"D5A101004E9E36C5CAF8A5F16B954891889D88AC88A0C8E040EAC8E5990DA94D",
            INIT_RAM_1D => X"2C95C6FB9F20CE3960D666B747CFA9A19329B8596FFEE1E024B142B177F2F304",
            INIT_RAM_1E => X"DE707BBF9C5F9F2C94F74F3878A3C0E77F38BF3CCB382E1A208EE6E77D77777C",
            INIT_RAM_1F => X"CFD000000FF1FDEA48C3E533DA331D77EE2A518E6F78B9C3B5CC2DD2EB3CED15",
            INIT_RAM_20 => X"352B1CB3ED3A7F8C2FFD607FCEBA3F08C9D6746F5995FADCAED4F9925B3995F3",
            INIT_RAM_21 => X"C99B2C66750F20C70263BBD92582182A4D582F00616B7CFB38D96C58229BA0F3",
            INIT_RAM_22 => X"9FE7EF999F9A613E9F3B221ADCF6DDED98B76C0411359EB7EA8B6CF7FD74DB39",
            INIT_RAM_23 => X"7FCC43F9E07FF5F7B7FFB7F43FFBAB30227FBFFADFCC229BB766E1E9BB1DD337",
            INIT_RAM_24 => X"F753B7D69DE33F40062F7CC2200006AB54007F9EFDFBFF36BBBB7D3F279EBD37",
            INIT_RAM_25 => X"53C5E2F714311FB17545D584A389DA684BD6EEC7C9727E7B3383FC3D9EA7FEEF",
            INIT_RAM_26 => X"9ABA0C567FB4EB3DDEEA2A35AA63453EE1ECF5A7F61F97F66CFD87E5F67B3F3E",
            INIT_RAM_27 => X"D17C7A32961E7478DFC018140683F37BFBFE7B72F66F6EFE9C173B3FFEF7ED26",
            INIT_RAM_28 => X"7AF88E7C0CFBEFB882E95651804688924D3403F93FED6BEF65D01BA62041FFF1",
            INIT_RAM_29 => X"C9178E5C66D2F7FFFFFCFEE7E9FBFFFFC0000002BFFFE3423CD538DC37AF239B",
            INIT_RAM_2A => X"41FD2ECFE6CD1FDBD37CEAE4EFCF5FD29B632B8FEFDE5C134AAADBB93D7CCE2C",
            INIT_RAM_2B => X"869FDDFB26DD2412BF6E5F332F3A3CF9FB9DA5E93C9FFEF6790F9E4EBFEFF7FC",
            INIT_RAM_2C => X"A3798FDB7FEB7A2ADA4B32ECFFE6AA889246099F76419D7208D39D7713DDA699",
            INIT_RAM_2D => X"526CB3DE4D9E4C9CB7F043828BC9F0AFDF2B7D5579BC7955454481DFF96EF8F0",
            INIT_RAM_2E => X"567B11080E43A75DC2158002801726EF841D647A75EF4449DD9B4696BE56749B",
            INIT_RAM_2F => X"DE014005764D523AEB374EA6D9B93FBAEB7A577E79C550E12F77762F3BF3DE09",
            INIT_RAM_30 => X"7757C5EF5492545AF576FEF75D9547FB1CD1CC50466056E8FE21E4FFF957CAC2",
            INIT_RAM_31 => X"5ADAD9E7CD3679F34D9A6CD379FBF26FCFD34EBAF4D3AEBFB2B2F795D5F5DFAB",
            INIT_RAM_32 => X"C357AC5224E91FBDDDAE6B91DCECD2668B1AFDFFFEEF7F4F7771524947BF65B2",
            INIT_RAM_33 => X"D0CBD11A22D0918161E9EFBA475FEEF342EFF7DDEFE7DFE9458C4FBF5BBE2E42",
            INIT_RAM_34 => X"DF7FAC98E34D5BAA0CD72E07DC6327FFDED8038DFFD8C9FFCC42E02BBE5EBE58",
            INIT_RAM_35 => X"89A70D55A17318A78ADD8BEF925534BC63257FB0D93EBF26FFAFAFD64F58CEDB",
            INIT_RAM_36 => X"674DD6BF7772BBFB7271F17BF7E9F0D04A728DC32DBD3A51CB83C8CECC468AEE",
            INIT_RAM_37 => X"EBF4D5555687F564A6BD5AE5FF3CB3F1E7F8EB559FCAA93B5236356090155131",
            INIT_RAM_38 => X"4132D95333C70B6F7E97BAD1336E66964FF55131FA52BB34E7D3FF91738E9DA8",
            INIT_RAM_39 => X"CF9A6CF3FD3FC6569BA7CFDECF3D1ACED3C7A3C7FBE7F6F3DDE1A9CF8DBADA3D",
            INIT_RAM_3A => X"F9E1EBDFC9FE79D006BEFC5EDE3FFF82FB4B22FA4DE351F4D3AEB9A6CF3E69B3",
            INIT_RAM_3B => X"AE555BD5B0D2D717BD367B0D9EEAB6ACF9FD1E95AC97F23B31BFF2774B31BA1F",
            INIT_RAM_3C => X"D5A101004E9E36C5CAF8A5F16B954891889D88AC88A0C8E040EAC8E5990DA94D",
            INIT_RAM_3D => X"2C95C6FB9F20CE3960D666B747CFA9A19329B8596FFEE1E024B142B177F2F304",
            INIT_RAM_3E => X"DE707BBF9C5F9F2C94F74F3878A3C0E77F38BF3CCB382E1A208EE6E77D77777C",
            INIT_RAM_3F => X"CFD000000FF1FDEA48C3E533DA331D77EE2A518E6F78B9C3B5CC2DD2EB3CED15"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"352B1CB3ED3A7F8C2FFD607FCEBA3F08C9D6746F5995FADCAED4F9925B3995F3",
            INIT_RAM_01 => X"C99B2C66750F20C70263BBD92582182A4D582F00616B7CFB38D96C58229BA0F3",
            INIT_RAM_02 => X"9FE7EF999F9A613E9F3B221ADCF6DDED98B76C0411359EB7EA8B6CF7FD74DB39",
            INIT_RAM_03 => X"7FCC43F9E07FF5F7B7FFB7F43FFBAB30227FBFFADFCC229BB766E1E9BB1DD337",
            INIT_RAM_04 => X"F753B7D69DE33F40062F7CC2200006AB54007F9EFDFBFF36BBBB7D3F279EBD37",
            INIT_RAM_05 => X"53C5E2F714311FB17545D584A389DA684BD6EEC7C9727E7B3383FC3D9EA7FEEF",
            INIT_RAM_06 => X"9ABA0C567FB4EB3DDEEA2A35AA63453EE1ECF5A7F61F97F66CFD87E5F67B3F3E",
            INIT_RAM_07 => X"D17C7A32961E7478DFC018140683F37BFBFE7B72F66F6EFE9C173B3FFEF7ED26",
            INIT_RAM_08 => X"7AF88E7C0CFBEFB882E95651804688924D3403F93FED6BEF65D01BA62041FFF1",
            INIT_RAM_09 => X"C9178E5C66D2F7FFFFFCFEE7E9FBFFFFC0000002BFFFE3423CD538DC37AF239B",
            INIT_RAM_0A => X"41FD2ECFE6CD1FDBD37CEAE4EFCF5FD29B632B8FEFDE5C134AAADBB93D7CCE2C",
            INIT_RAM_0B => X"869FDDFB26DD2412BF6E5F332F3A3CF9FB9DA5E93C9FFEF6790F9E4EBFEFF7FC",
            INIT_RAM_0C => X"A3798FDB7FEB7A2ADA4B32ECFFE6AA889246099F76419D7208D39D7713DDA699",
            INIT_RAM_0D => X"526CB3DE4D9E4C9CB7F043828BC9F0AFDF2B7D5579BC7955454481DFF96EF8F0",
            INIT_RAM_0E => X"567B11080E43A75DC2158002801726EF841D647A75EF4449DD9B4696BE56749B",
            INIT_RAM_0F => X"DE014005764D523AEB374EA6D9B93FBAEB7A577E79C550E12F77762F3BF3DE09",
            INIT_RAM_10 => X"7757C5EF5492545AF576FEF75D9547FB1CD1CC50466056E8FE21E4FFF957CAC2",
            INIT_RAM_11 => X"5ADAD9E7CD3679F34D9A6CD379FBF26FCFD34EBAF4D3AEBFB2B2F795D5F5DFAB",
            INIT_RAM_12 => X"C357AC5224E91FBDDDAE6B91DCECD2668B1AFDFFFEEF7F4F7771524947BF65B2",
            INIT_RAM_13 => X"D0CBD11A22D0918161E9EFBA475FEEF342EFF7DDEFE7DFE9458C4FBF5BBE2E42",
            INIT_RAM_14 => X"DF7FAC98E34D5BAA0CD72E07DC6327FFDED8038DFFD8C9FFCC42E02BBE5EBE58",
            INIT_RAM_15 => X"89A70D55A17318A78ADD8BEF925534BC63257FB0D93EBF26FFAFAFD64F58CEDB",
            INIT_RAM_16 => X"674DD6BF7772BBFB7271F17BF7E9F0D04A728DC32DBD3A51CB83C8CECC468AEE",
            INIT_RAM_17 => X"EBF4D5555687F564A6BD5AE5FF3CB3F1E7F8EB559FCAA93B5236356090155131",
            INIT_RAM_18 => X"4132D95333C70B6F7E97BAD1336E66964FF55131FA52BB34E7D3FF91738E9DA8",
            INIT_RAM_19 => X"CF9A6CF3FD3FC6569BA7CFDECF3D1ACED3C7A3C7FBE7F6F3DDE1A9CF8DBADA3D",
            INIT_RAM_1A => X"F9E1EBDFC9FE79D006BEFC5EDE3FFF82FB4B22FA4DE351F4D3AEB9A6CF3E69B3",
            INIT_RAM_1B => X"AE555BD5B0D2D717BD367B0D9EEAB6ACF9FD1E95AC97F23B31BFF2774B31BA1F",
            INIT_RAM_1C => X"D5A101004E9E36C5CAF8A5F16B954891889D88AC88A0C8E040EAC8E5990DA94D",
            INIT_RAM_1D => X"2C95C6FB9F20CE3960D666B747CFA9A19329B8596FFEE1E024B142B177F2F304",
            INIT_RAM_1E => X"DE707BBF9C5F9F2C94F74F3878A3C0E77F38BF3CCB382E1A208EE6E77D77777C",
            INIT_RAM_1F => X"CFD000000FF1FDEA48C3E533DA331D77EE2A518E6F78B9C3B5CC2DD2EB3CED15",
            INIT_RAM_20 => X"352B1CB3ED3A7F8C2FFD607FCEBA3F08C9D6746F5995FADCAED4F9925B3995F3",
            INIT_RAM_21 => X"C99B2C66750F20C70263BBD92582182A4D582F00616B7CFB38D96C58229BA0F3",
            INIT_RAM_22 => X"9FE7EF999F9A613E9F3B221ADCF6DDED98B76C0411359EB7EA8B6CF7FD74DB39",
            INIT_RAM_23 => X"7FCC43F9E07FF5F7B7FFB7F43FFBAB30227FBFFADFCC229BB766E1E9BB1DD337",
            INIT_RAM_24 => X"F753B7D69DE33F40062F7CC2200006AB54007F9EFDFBFF36BBBB7D3F279EBD37",
            INIT_RAM_25 => X"53C5E2F714311FB17545D584A389DA684BD6EEC7C9727E7B3383FC3D9EA7FEEF",
            INIT_RAM_26 => X"9ABA0C567FB4EB3DDEEA2A35AA63453EE1ECF5A7F61F97F66CFD87E5F67B3F3E",
            INIT_RAM_27 => X"D17C7A32961E7478DFC018140683F37BFBFE7B72F66F6EFE9C173B3FFEF7ED26",
            INIT_RAM_28 => X"7AF88E7C0CFBEFB882E95651804688924D3403F93FED6BEF65D01BA62041FFF1",
            INIT_RAM_29 => X"C9178E5C66D2F7FFFFFCFEE7E9FBFFFFC0000002BFFFE3423CD538DC37AF239B",
            INIT_RAM_2A => X"41FD2ECFE6CD1FDBD37CEAE4EFCF5FD29B632B8FEFDE5C134AAADBB93D7CCE2C",
            INIT_RAM_2B => X"869FDDFB26DD2412BF6E5F332F3A3CF9FB9DA5E93C9FFEF6790F9E4EBFEFF7FC",
            INIT_RAM_2C => X"A3798FDB7FEB7A2ADA4B32ECFFE6AA889246099F76419D7208D39D7713DDA699",
            INIT_RAM_2D => X"526CB3DE4D9E4C9CB7F043828BC9F0AFDF2B7D5579BC7955454481DFF96EF8F0",
            INIT_RAM_2E => X"567B11080E43A75DC2158002801726EF841D647A75EF4449DD9B4696BE56749B",
            INIT_RAM_2F => X"DE014005764D523AEB374EA6D9B93FBAEB7A577E79C550E12F77762F3BF3DE09",
            INIT_RAM_30 => X"7757C5EF5492545AF576FEF75D9547FB1CD1CC50466056E8FE21E4FFF957CAC2",
            INIT_RAM_31 => X"5ADAD9E7CD3679F34D9A6CD379FBF26FCFD34EBAF4D3AEBFB2B2F795D5F5DFAB",
            INIT_RAM_32 => X"C357AC5224E91FBDDDAE6B91DCECD2668B1AFDFFFEEF7F4F7771524947BF65B2",
            INIT_RAM_33 => X"D0CBD11A22D0918161E9EFBA475FEEF342EFF7DDEFE7DFE9458C4FBF5BBE2E42",
            INIT_RAM_34 => X"DF7FAC98E34D5BAA0CD72E07DC6327FFDED8038DFFD8C9FFCC42E02BBE5EBE58",
            INIT_RAM_35 => X"89A70D55A17318A78ADD8BEF925534BC63257FB0D93EBF26FFAFAFD64F58CEDB",
            INIT_RAM_36 => X"674DD6BF7772BBFB7271F17BF7E9F0D04A728DC32DBD3A51CB83C8CECC468AEE",
            INIT_RAM_37 => X"EBF4D5555687F564A6BD5AE5FF3CB3F1E7F8EB559FCAA93B5236356090155131",
            INIT_RAM_38 => X"4132D95333C70B6F7E97BAD1336E66964FF55131FA52BB34E7D3FF91738E9DA8",
            INIT_RAM_39 => X"CF9A6CF3FD3FC6569BA7CFDECF3D1ACED3C7A3C7FBE7F6F3DDE1A9CF8DBADA3D",
            INIT_RAM_3A => X"F9E1EBDFC9FE79D006BEFC5EDE3FFF82FB4B22FA4DE351F4D3AEB9A6CF3E69B3",
            INIT_RAM_3B => X"AE555BD5B0D2D717BD367B0D9EEAB6ACF9FD1E95AC97F23B31BFF2774B31BA1F",
            INIT_RAM_3C => X"D5A101004E9E36C5CAF8A5F16B954891889D88AC88A0C8E040EAC8E5990DA94D",
            INIT_RAM_3D => X"2C95C6FB9F20CE3960D666B747CFA9A19329B8596FFEE1E024B142B177F2F304",
            INIT_RAM_3E => X"DE707BBF9C5F9F2C94F74F3878A3C0E77F38BF3CCB382E1A208EE6E77D77777C",
            INIT_RAM_3F => X"CFD000000FF1FDEA48C3E533DA331D77EE2A518E6F78B9C3B5CC2DD2EB3CED15"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"1DC552A39BB3FC75E7D79B3AC5FF29E6FF24FDCECEF9FFB3B31D9B090909075F",
            INIT_RAM_01 => X"A6512ADBE8C8610EDB9DCDC020CD6E58E6DAA2A3B64FA4BBDE0BE5D3DF269ACF",
            INIT_RAM_02 => X"64D432F9D8FAEBA58FCF1478652846717F596FB523EE6BF9EB2E935B5D942424",
            INIT_RAM_03 => X"BBD276BCB925DA281B2C6E6CF3ACC893C0419D721A34C2DCEF1AEDE6777F9971",
            INIT_RAM_04 => X"D14B49CAE29B565578B64AE94AA5BEBED0104DF69D7577FCB557CF696B5F54DC",
            INIT_RAM_05 => X"8BA53D5545AD27F087F3F0544E5EA5B780BC6B1BA32DB44F44D598B728A68C53",
            INIT_RAM_06 => X"553BBFBA1764200E04FA9E64D1D2F70A3EE7264508A3E3931BD9367E15D2CDF7",
            INIT_RAM_07 => X"482F9B95A99B77F7E375B0D603BD3020FA83FD5BBC7E375B0D423E186CF0BE1C",
            INIT_RAM_08 => X"7FF5CF1530E1E3DECE86E2A9A4C22412980781C08544E90010F863B49F4447C4",
            INIT_RAM_09 => X"F3BFF8F5F5D7E2B2A2BB3ABF9FE5A5E99D5D3BBD6DF735F47FFB7E49F6FF6CDF",
            INIT_RAM_0A => X"4CC4A99B9033A2795A1FDEE8EFC67AC373F37D7593FCCF45ACDA11A24B7BF2B0",
            INIT_RAM_0B => X"B721A234B170B967B967C97EFF2F967D6B72C6B61E21FD74CC2E0034FEF994AE",
            INIT_RAM_0C => X"9E7FFE13F21DFDA43EEC33C2E1F370F9FEEF619DFFFFF132865FE7CD5FACCDDC",
            INIT_RAM_0D => X"C7DB0C04142BB77E4BFCFB37FAE76DD3F25AFF9FCBDCE1EC9D3CBD74C4A7CFDB",
            INIT_RAM_0E => X"818EAA7FAC81A79C67EC364440D6FFFFF9D86434D7DEA14599F64E1BC0004C49",
            INIT_RAM_0F => X"11DB36B5C97D836F3E33E3EAA19F2D7B26E27A4C1130DC6D6D6F6D6F6F6CAFFA",
            INIT_RAM_10 => X"003EEBAE8151BB843E1ED3CA74E27A4C1171BAE91D9A431B7B5C97E0DB6FF245",
            INIT_RAM_11 => X"9A366E98058A1866C85B3E7F9CF1BFFE79E34514111110405505115544011441",
            INIT_RAM_12 => X"FAE7D7975CEF0F7AAE95944AF29C59CD086C2BBF353FE1230D86C3719B6D95AD",
            INIT_RAM_13 => X"24A45EFD22E4218E777E61F1337FE736AADA688C0E5BB57E9DBB7F7DF757D6AE",
            INIT_RAM_14 => X"427B66A21704C7B3DB30A8098A80D42A3CCABA847B96D73B7A9D6D18E63508BF",
            INIT_RAM_15 => X"EA8882576A3BB0D3825C802FEBF5CAACCF69F5259B993A8E1495FE90B93D47B7",
            INIT_RAM_16 => X"BF80C05B3E4C4AE798631FD67CD5CBB94D66759C35E2AF692968B0515B57397E",
            INIT_RAM_17 => X"153B14B91EC14657857BED800920001FCC7E9A4ED039A618C1A4CC241348F35F",
            INIT_RAM_18 => X"77BBB0E8567A1598A85605CEB74B92ABABA2823F4090505E95100D4BCFE8C3E2",
            INIT_RAM_19 => X"CA873DC485292E948251DF549A44C775D35E879D9C01299C2693B0F8DE766736",
            INIT_RAM_1A => X"A36370B752D18367871942F11BD275E45FC3F977DF5EFCF9E8C0E57F4F32732E",
            INIT_RAM_1B => X"FF63323F35B72F6DBDBFF6CC4A40884BA8846E69E6D584D84DFDFB9368D6B7AD",
            INIT_RAM_1C => X"6E7F6F377ECFACBA7F6BADF752E51FA7FF9258FF9ABBFFCCDFFFFE6FFDF91F98",
            INIT_RAM_1D => X"D24BB73ACCD6726F4E99ABAFA69E7BBA99A4D2D7392667D674A774CFFD936FB7",
            INIT_RAM_1E => X"E7FFE6A35DFC849247A5735645524D24BCEB335E73337860CD04924335645524",
            INIT_RAM_1F => X"EA38FBF08D3F7C2C9A7AEBCBBA99A734F7774DD2DB67F4DCFECFF4D81C6BBF9C",
            INIT_RAM_20 => X"E33C5FFB7F93A73F3CFFAFFDD766CD2EBB3669F7E7EA6B2109C209F1C2047389",
            INIT_RAM_21 => X"D5F1EDBB963ACEDC7D987CCB735C5BFDD42C9FDCD738FFC64FFFF801797E77D9",
            INIT_RAM_22 => X"02EA1911D90011A5750B3F0A48EABD5BB2BFCB66AFDD545BB4ADAF3BDCBD4765",
            INIT_RAM_23 => X"F80F800C1CF84DEEDEE74E2D1E7DBF7B79F3F934CABEEFCFFDFBD2584E4C0309",
            INIT_RAM_24 => X"AC684A74A9B04F6A148152C8925097B50D34FCA727E7C88888888DFEBEF9415C",
            INIT_RAM_25 => X"1400158B2CFBDB32AE28ACFBCD45009FF557488F62BED53691800077674D05BC",
            INIT_RAM_26 => X"9FF33C5F204AE65ADE6710B203AB175BAAFBD639567DBC196FDDA011BAA40097",
            INIT_RAM_27 => X"4DA71155BACCC148DAD786B205392CAF056FC2B2A021D15F98476DEE15E415D2",
            INIT_RAM_28 => X"AC774BA4E001EC16C9817947A2065565A2B2917608A2F912FE93ED82BEC7E71C",
            INIT_RAM_29 => X"DB2DB13B52DBE67EF6FA05F33F769A05DEE1A6368A92C9DAD9F55D6D5D88EAFB",
            INIT_RAM_2A => X"D77EF96D9EDDFF3737B6CB9B9FDA8ED436E9726B73E6DBFC91DCD9BA0FB3A89C",
            INIT_RAM_2B => X"27027DB3B679286FD5FECEFDADA4CBED0983CFDE9E56F1B0DAC3ED7A78C38F3F",
            INIT_RAM_2C => X"77CCECE01581F777C17A68CC08C9164BA164BAFE8B327A81E64E71823A81AE50",
            INIT_RAM_2D => X"99911F011E266444D312309C3445FD3E371DF544449CCD75B5675EA9E96F60C7",
            INIT_RAM_2E => X"00007E48DEFC7B2CD1F4DD550DCE6737463504448A18E9115BE535B4EE42B050",
            INIT_RAM_2F => X"5ED9B8378E1DCDE392CE6732FC28DF29F1F3DDA827B44F672BCFE56C0CCC8000",
            INIT_RAM_30 => X"4ED5DE57D641E0FD979F80701936BABB7426E580E1B6E3266DD0C7724CF6BBCA",
            INIT_RAM_31 => X"D574B3719E1A5ECF54DCBDD5AF14A31B17F1C92DD5970256FABF5EA9F974DC57",
            INIT_RAM_32 => X"15BC0CB69FACB2CB4EF9B700A78A3CF735CA9FDF7AE19BE151E5FDE67EEE67F0",
            INIT_RAM_33 => X"1EFFF0B22D0021DD0AE970A5419180808EFA4D48BE46472761B7B3E96E4B55C5",
            INIT_RAM_34 => X"D1F48F58D1EB9561A27C32A1947FD7F61DF75D64ABFF43640689FF2100C7214B",
            INIT_RAM_35 => X"10610236B76C5B16FDED44FBCCDFA46A0F76B17312FBF05CAF23610485426D84",
            INIT_RAM_36 => X"6FFDBDA6B143DFE9FFBA9FBC3110B08BDB55C3023E77FDEFF32BFF72BFFB2BF9",
            INIT_RAM_37 => X"67B0EFB800C9FFBC6AFBB6D9CE7AB39267DDBE56F64E79C4E957A6FDDFBE5F7D",
            INIT_RAM_38 => X"EBF5DEDCE8CCB5F5A2FE754772E49DB479FEFA605ED4B7F1E4184D3E38A003FE",
            INIT_RAM_39 => X"FE7F2CD7FCBFDC7FE7D49D5EAB3F381FDB8F5E05ADA889F9F11000780FDF7A77",
            INIT_RAM_3A => X"70E9C37CBB6EB6E4F6D793D6BBBB699DA21018A3D03448693833EF3D650FD65E",
            INIT_RAM_3B => X"4D2C33E926EAE9D5D7F9DDDBE8EEDCD6654E47B16FBD126023C19AE37DE5D3CE",
            INIT_RAM_3C => X"75A857EE1171F8EB578C6FDD8C58E6EB03BB1816B949950F8423B986B6D6D6D2",
            INIT_RAM_3D => X"855C7D42726EBCA691146A85AF5C46C6760EB71C730FEBF719E6EE3EEDD70D6B",
            INIT_RAM_3E => X"75E52F2166F040B063E081039FF784CB060314224C14934541307A40277FB1C9",
            INIT_RAM_3F => X"B4C97E5FF22AF024CB00880088009ED9788D32B7EB47BB9F8AB9FBC7BCC1E133"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_2,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"4845BD5B243DAED2B2489B313A35C50252AFD0FFB76FE7342335FFF132FD92FF",
            INIT_RAM_01 => X"5372B72B484E2F2664B735B69A5AB532B086BA4C62AD6D56EECBDB6984B25145",
            INIT_RAM_02 => X"DD6E630C15271E48CA801988654FB501D5393392EE765C1EC95C1E4D86F18A96",
            INIT_RAM_03 => X"17F7F5724D40707E6FF30002982023020449B4680C45D1CFAD8EB30A061DB8FE",
            INIT_RAM_04 => X"BD52921D249E377EDBD14EA309EEDAA57DA85F55DBB7048A69A4C801013948B6",
            INIT_RAM_05 => X"5E2B1A3E16869E1D37BCE906B82F401CBD467617DB34D9E0C80B5E6E10063EC4",
            INIT_RAM_06 => X"BA611013110188547995B108BB2DAE76F4A3A0D98845F9248BDFA45E10CA403A",
            INIT_RAM_07 => X"D0734B461A36980411EB2A6C1BE76029258777EF227A8F6E84F74C4436098F67",
            INIT_RAM_08 => X"60A229B98541E6FE734DE2280A9B57FCD5A9BEFEF7CDA5ABEB44FD73D2794D56",
            INIT_RAM_09 => X"84735325ACC969B2EAE10A1478D866FA67DDEF7BBF75E6958B6D02DC6D0F8076",
            INIT_RAM_0A => X"7833830C7B2C7AFB8A8D203C312306DA0E72641FFB93D79B5EC04F44AD55F4B8",
            INIT_RAM_0B => X"1C387A7970C7F3E688673CF5975EE3E5FF105CFCCF9F725D698FB088B063063C",
            INIT_RAM_0C => X"96CE81973CB55590446D599375501366EC343561BCF83357F8823671393B278C",
            INIT_RAM_0D => X"8CEBCB187AE5D44ECA689C9BD4E5AE544DEA7E90D186B9F335F3223877AAD541",
            INIT_RAM_0E => X"BCCF19EEF299751C919C9C13C6FB9ED711AC4DA7D947CC79E9B6323EF6CE6263",
            INIT_RAM_0F => X"763DD7AAFEED3F4AD4EA7491ADE6F14E6DBADD0F090A8DF34D7BAD35DD2275F0",
            INIT_RAM_10 => X"37309C08305A10187707E3D57DDE4931F1D9E97A8F378981ABBF8D7B6B7549C3",
            INIT_RAM_11 => X"9467DA6C480E6D19CEEA8451CEFA88FD70E7925B0302F877F87FA833FBD147E9",
            INIT_RAM_12 => X"99716B8CBAE953D061FAC3D6337D5BA4D6D7090929944AB6FA3357801066B658",
            INIT_RAM_13 => X"F331598B364EF27516CC49A4662C5E5C92ED140D96372E7A7833AE4346982375",
            INIT_RAM_14 => X"A5875745B625C6CA7A7292332492D139728A689DA1AE78B6B44CE4F4A4EA5A22",
            INIT_RAM_15 => X"CD2E1AF14C30545297A91BED3AEAEFF8F696B5F4FC80BC6B1A2559492E9198E4",
            INIT_RAM_16 => X"75B74FB9AF7C1A492952F7EEAA0E7CF9FBEDD0FB47EEFDCC3734B816F355C913",
            INIT_RAM_17 => X"88537A811D4EF6CD9668CCD3E2E7A8041788DCA5F7E08AF52AF527607BF06DEB",
            INIT_RAM_18 => X"66591A35ADD26B6B7E33CA56E9A4759EFA7E68F98AE7CE9507755C74C430286A",
            INIT_RAM_19 => X"56F9FDFE7D64C1F4E1F5641845CD17E836B97780400C702723FA8E7C7BBD6F06",
            INIT_RAM_1A => X"0A01FDC7FE2CBF038A61DEA5FCE2C10C8F35FBF80C05ABFF4B6935287B125E8D",
            INIT_RAM_1B => X"607D53A5C955D5D1412F8361617A5444E971FD187442A60FB04457857BECC312",
            INIT_RAM_1C => X"CE4B65409D6F079D709A56C38DC3BCEF07459A416EB4E8F3D73CC714F4333AFE",
            INIT_RAM_1D => X"04B57D8E0D755851232838F9B5348838530D7AF95411555D263B8CA86A5D29D7",
            INIT_RAM_1E => X"DF7D7BF31C6072BFA7993996AB7DD2F3EE4009844CC9D6CF9E583AEC48A52F29",
            INIT_RAM_1F => X"1EEA3633EFEA856D05BA968C1B3C30CA1788DD95D16B8F914DDDFC3EE5C69945",
            INIT_RAM_20 => X"95DE707778B17C2379847A23AE6B8BB01F36F3F44A8162566D9FB15DE7CC83F7",
            INIT_RAM_21 => X"EEC890579E95D5A0A546CCCDD48577558ABE7CA36EF67A70F6A8758BDA052D5B",
            INIT_RAM_22 => X"6BAD12FDFB527EF4F87F4A23EC13CBC0262D8899A3A290F04F41C1324045B9FC",
            INIT_RAM_23 => X"85287860729C77B6C68CAEA3033A6E84D67249B594C407B39C68B4C1C97FDEFC",
            INIT_RAM_24 => X"CB76FAB179E9619BC7E7E9C9FD801CF87DBA1EA496E829D4E62861E1AF436A75",
            INIT_RAM_25 => X"65F627A15E1057ADEE7B9E27122A58FF2B98B1EA560390C7E8F715861814E04D",
            INIT_RAM_26 => X"0004406BD60A023AB063D4E5966EA41AA997F5A49BFCB1657A9732D28EB8217E",
            INIT_RAM_27 => X"4ED4AE2B1650D21EAFE01E7099EFCA3094FD4D705CF6B84AE21583E13385F865",
            INIT_RAM_28 => X"5725EA43CE18F187A1DE4DAABEA97963E3A7A96B8B7CBC095BEB7CE46274D9AF",
            INIT_RAM_29 => X"3C563C8B02C8CC39C64DDCEA1BEEB5E7353F93786145598FE634EF1000179B34",
            INIT_RAM_2A => X"735AF87DAE59FABBD7DEAF8717F2B72F428F5E37E5D6E13157B99CBD2D73B9C7",
            INIT_RAM_2B => X"9555AFBBD3AEBFCABFBBED7A5C5FE9BD0E6A91C6E7610042695EEB08D8881B1D",
            INIT_RAM_2C => X"C5595549AC64787878F5CE14C664CF9EB0CDAFFBABEF1E83358371B9ED96E506",
            INIT_RAM_2D => X"CAE30B9FE6AA29FFF6F72DA73DFE4F7ACD39687B9E69C5359E9B991F0746EFFB",
            INIT_RAM_2E => X"EFEF92C2FA4D8D4E4AC86C277338FA37BCDD9D47781EDBAF7FC03C1BCD23D0AF",
            INIT_RAM_2F => X"E629BDF93D7F5B5BAF92FBAB477E9B315DB5A310CFACC7408DF9A544B1E57AF6",
            INIT_RAM_30 => X"3F1BF746FBFFC353E37263FF38A796EF39E3FD7DFEBA7FFEFFBF17ABAF09E909",
            INIT_RAM_31 => X"636CDEB4BDFCAEEFC61DFFEFB7E26262DEF2CB9F71565824FEBF3F7BDDEABB59",
            INIT_RAM_32 => X"FF9FFF6E3881C81AFDCF2257FD4F8ED5257D0E9B800726B646C8A8E5012F76DF",
            INIT_RAM_33 => X"4E93FD3C1238FFAFBD7FDF567FA8FEF024F33AFD3AABC6B105EA80272D64895F",
            INIT_RAM_34 => X"47B2AFF5B87AA26AFFDD317DEDCFBDFFE1A0CAD3B58877DD2F647F7DF748E7CF",
            INIT_RAM_35 => X"6F6DFFF29CB70FFD25A59DFFFED7B3F7E8B4CE6FFF3EF9CEC6BAE57ABFFFCEE6",
            INIT_RAM_36 => X"AEC4837C2A5FECBB94C1C969FFDDFF79BFFAAFDCA8D748399ABF75558ADD02F5",
            INIT_RAM_37 => X"DDE6FC8EBE3F9F3C3DFC6E8F07BFD31D50660B1E0B2506A533CE0E340C7C745C",
            INIT_RAM_38 => X"8E33E171D3C17C17D665B4DC7E31C7957667EB9A44CE0EEDBBBD391D3128AAA3",
            INIT_RAM_39 => X"8CE19D963783FC4F1D83AC65DFF0E6661186734DB8C4580E23E97CDCD8FF66DD",
            INIT_RAM_3A => X"A8AE5EF365D000000C86C7866B1BF5398C30634E3D04A901DF994261B3D4BEFF",
            INIT_RAM_3B => X"80000000F3379EE5ADE3DD0111DC4D877F2C1BE8E59CF7F73AA8D565B9B6FAA5",
            INIT_RAM_3C => X"000000000000000000000000001ED5A9AB3575A6DFE371D6AFE4F82C6516249B",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"8000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"3C00000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"97B6A1C61A005A50A952155B13C5545DD3BEC93BE9D969D8A0ECD699493B0999",
            INIT_RAM_01 => X"3662D18D53B5529C6B462D904030410F2987F76AE99082301A76DFFCDBD280F8",
            INIT_RAM_02 => X"B9C0D70012C8100F02A57E94F585103548FF1A788E13666C0FB4D30C24833694",
            INIT_RAM_03 => X"A5449038F03B7FEE480307F1102CC52451C0C25B0829B0EEFDE03D3D04142A51",
            INIT_RAM_04 => X"1854A05040027D0002B7F59B59C74C1766AA3151C10A1F5823656671E023EDE4",
            INIT_RAM_05 => X"F1D0AF734000640F8BAD82B5BAA3880AC05C0BDC7B96FE9AF64C00BA23C80332",
            INIT_RAM_06 => X"8324E2621D8F4B2578AEE658FF1EA65185D11F0800600588B1001801688C402E",
            INIT_RAM_07 => X"DA0F9D292022728848197B2E8F96145887303588887D43171EA08207E2C32C08",
            INIT_RAM_08 => X"A3D5A2576AABAEBBA1EA5AE10DAAD52414511401400DADA8096002B29A3DD539",
            INIT_RAM_09 => X"3726B597AA78A800C841394877FBFFFFFFEFFFEA95559D4C16AFD65F97EA7A28",
            INIT_RAM_0A => X"6A1347C1D90061090065BFF375FDD0F8E988E4274031B1887FC3E66678809F45",
            INIT_RAM_0B => X"000F6677ACE21AC02FE7209AEDA8CB4201B4F1766126054967611195182E7D90",
            INIT_RAM_0C => X"8D662F3EC87ED1491AF32277F3C0BB100148622E0CDF73EACE41E12A61721B80",
            INIT_RAM_0D => X"A99736C201F09D0F807491FC11C7647DDB62BB24B293E68999B65D7081DF3252",
            INIT_RAM_0E => X"808272F5F5A954A45BB83A775740002AC682D4010C5355C23772E82D0FA87E35",
            INIT_RAM_0F => X"29AE35540024894036BD6D5B6A48126C0254A5FC845007121155575652C0B774",
            INIT_RAM_10 => X"62280010246122210C8D050D801929C3A10032DADD79E0AD0A48282D89E28C59",
            INIT_RAM_11 => X"10A8A09916C82645B26C932582440590706C92449B24912012A008075E01882C",
            INIT_RAM_12 => X"F1F78129454A607B0294BDE97ED3640C5746110020B09020826699949A044181",
            INIT_RAM_13 => X"474C99DFB9715D37CF22B3EB29400C45E5000C161250A040225662BF02FE98D6",
            INIT_RAM_14 => X"2016DB528401BC1B31089935A880991602031CB2016C32040CDF193E8200488A",
            INIT_RAM_15 => X"C9BE7DDDCEC45069CCBE50C429BE506ECA3FAA156040A204D942536D920008DD",
            INIT_RAM_16 => X"962428A4C940CFFAC08EA2852A2A25AB0C80525581438E71F62A61D3BF72059B",
            INIT_RAM_17 => X"4A40195556EFFC488C732D5A852224C889B340095CBC508A4199066D714D34A8",
            INIT_RAM_18 => X"8CC93C708006AC721B862318602C01212258D2CE44080C0911B7FFE488384011",
            INIT_RAM_19 => X"1664B20582486B096DC93F761554AC21ED5A1832824B345B423A3401565022D3",
            INIT_RAM_1A => X"E39A83371278E663BC0B1BF1E5E1000D2436C540240078096C03664B205992C8",
            INIT_RAM_1B => X"25311085A8A28353CC9EC427B10012FCB7ECF51905B4349160D5C48CB20EA029",
            INIT_RAM_1C => X"422B02856A0C0AD1CA3495D96324C224420C4208C200C2A15962E86D50CD21FC",
            INIT_RAM_1D => X"F056013D840BAFC5BD89015A00028449C55865048F8D12B483CCB84C224D8C69",
            INIT_RAM_1E => X"5AD625192CA1B0B2EF37EA310192F34A325946F20F4CD1DBB456EE63C1999820",
            INIT_RAM_1F => X"52D00000019FE208805BFE601398005F7A9801BFFFFBFF730FFE51772412ED29",
            INIT_RAM_20 => X"97B6A1C61A005A50A952155B13C5545DD3BEC93BE9D969D8A0ECD699493B0999",
            INIT_RAM_21 => X"3662D18D53B5529C6B462D904030410F2987F76AE99082301A76DFFCDBD280F8",
            INIT_RAM_22 => X"B9C0D70012C8100F02A57E94F585103548FF1A788E13666C0FB4D30C24833694",
            INIT_RAM_23 => X"A5449038F03B7FEE480307F1102CC52451C0C25B0829B0EEFDE03D3D04142A51",
            INIT_RAM_24 => X"1854A05040027D0002B7F59B59C74C1766AA3151C10A1F5823656671E023EDE4",
            INIT_RAM_25 => X"F1D0AF734000640F8BAD82B5BAA3880AC05C0BDC7B96FE9AF64C00BA23C80332",
            INIT_RAM_26 => X"8324E2621D8F4B2578AEE658FF1EA65185D11F0800600588B1001801688C402E",
            INIT_RAM_27 => X"DA0F9D292022728848197B2E8F96145887303588887D43171EA08207E2C32C08",
            INIT_RAM_28 => X"A3D5A2576AABAEBBA1EA5AE10DAAD52414511401400DADA8096002B29A3DD539",
            INIT_RAM_29 => X"3726B597AA78A800C841394877FBFFFFFFEFFFEA95559D4C16AFD65F97EA7A28",
            INIT_RAM_2A => X"6A1347C1D90061090065BFF375FDD0F8E988E4274031B1887FC3E66678809F45",
            INIT_RAM_2B => X"000F6677ACE21AC02FE7209AEDA8CB4201B4F1766126054967611195182E7D90",
            INIT_RAM_2C => X"8D662F3EC87ED1491AF32277F3C0BB100148622E0CDF73EACE41E12A61721B80",
            INIT_RAM_2D => X"A99736C201F09D0F807491FC11C7647DDB62BB24B293E68999B65D7081DF3252",
            INIT_RAM_2E => X"808272F5F5A954A45BB83A775740002AC682D4010C5355C23772E82D0FA87E35",
            INIT_RAM_2F => X"29AE35540024894036BD6D5B6A48126C0254A5FC845007121155575652C0B774",
            INIT_RAM_30 => X"62280010246122210C8D050D801929C3A10032DADD79E0AD0A48282D89E28C59",
            INIT_RAM_31 => X"10A8A09916C82645B26C932582440590706C92449B24912012A008075E01882C",
            INIT_RAM_32 => X"F1F78129454A607B0294BDE97ED3640C5746110020B09020826699949A044181",
            INIT_RAM_33 => X"474C99DFB9715D37CF22B3EB29400C45E5000C161250A040225662BF02FE98D6",
            INIT_RAM_34 => X"2016DB528401BC1B31089935A880991602031CB2016C32040CDF193E8200488A",
            INIT_RAM_35 => X"C9BE7DDDCEC45069CCBE50C429BE506ECA3FAA156040A204D942536D920008DD",
            INIT_RAM_36 => X"962428A4C940CFFAC08EA2852A2A25AB0C80525581438E71F62A61D3BF72059B",
            INIT_RAM_37 => X"4A40195556EFFC488C732D5A852224C889B340095CBC508A4199066D714D34A8",
            INIT_RAM_38 => X"8CC93C708006AC721B862318602C01212258D2CE44080C0911B7FFE488384011",
            INIT_RAM_39 => X"1664B20582486B096DC93F761554AC21ED5A1832824B345B423A3401565022D3",
            INIT_RAM_3A => X"E39A83371278E663BC0B1BF1E5E1000D2436C540240078096C03664B205992C8",
            INIT_RAM_3B => X"25311085A8A28353CC9EC427B10012FCB7ECF51905B4349160D5C48CB20EA029",
            INIT_RAM_3C => X"422B02856A0C0AD1CA3495D96324C224420C4208C200C2A15962E86D50CD21FC",
            INIT_RAM_3D => X"F056013D840BAFC5BD89015A00028449C55865048F8D12B483CCB84C224D8C69",
            INIT_RAM_3E => X"5AD625192CA1B0B2EF37EA310192F34A325946F20F4CD1DBB456EE63C1999820",
            INIT_RAM_3F => X"52D00000019FE208805BFE601398005F7A9801BFFFFBFF730FFE51772412ED29"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"97B6A1C61A005A50A952155B13C5545DD3BEC93BE9D969D8A0ECD699493B0999",
            INIT_RAM_01 => X"3662D18D53B5529C6B462D904030410F2987F76AE99082301A76DFFCDBD280F8",
            INIT_RAM_02 => X"B9C0D70012C8100F02A57E94F585103548FF1A788E13666C0FB4D30C24833694",
            INIT_RAM_03 => X"A5449038F03B7FEE480307F1102CC52451C0C25B0829B0EEFDE03D3D04142A51",
            INIT_RAM_04 => X"1854A05040027D0002B7F59B59C74C1766AA3151C10A1F5823656671E023EDE4",
            INIT_RAM_05 => X"F1D0AF734000640F8BAD82B5BAA3880AC05C0BDC7B96FE9AF64C00BA23C80332",
            INIT_RAM_06 => X"8324E2621D8F4B2578AEE658FF1EA65185D11F0800600588B1001801688C402E",
            INIT_RAM_07 => X"DA0F9D292022728848197B2E8F96145887303588887D43171EA08207E2C32C08",
            INIT_RAM_08 => X"A3D5A2576AABAEBBA1EA5AE10DAAD52414511401400DADA8096002B29A3DD539",
            INIT_RAM_09 => X"3726B597AA78A800C841394877FBFFFFFFEFFFEA95559D4C16AFD65F97EA7A28",
            INIT_RAM_0A => X"6A1347C1D90061090065BFF375FDD0F8E988E4274031B1887FC3E66678809F45",
            INIT_RAM_0B => X"000F6677ACE21AC02FE7209AEDA8CB4201B4F1766126054967611195182E7D90",
            INIT_RAM_0C => X"8D662F3EC87ED1491AF32277F3C0BB100148622E0CDF73EACE41E12A61721B80",
            INIT_RAM_0D => X"A99736C201F09D0F807491FC11C7647DDB62BB24B293E68999B65D7081DF3252",
            INIT_RAM_0E => X"808272F5F5A954A45BB83A775740002AC682D4010C5355C23772E82D0FA87E35",
            INIT_RAM_0F => X"29AE35540024894036BD6D5B6A48126C0254A5FC845007121155575652C0B774",
            INIT_RAM_10 => X"62280010246122210C8D050D801929C3A10032DADD79E0AD0A48282D89E28C59",
            INIT_RAM_11 => X"10A8A09916C82645B26C932582440590706C92449B24912012A008075E01882C",
            INIT_RAM_12 => X"F1F78129454A607B0294BDE97ED3640C5746110020B09020826699949A044181",
            INIT_RAM_13 => X"474C99DFB9715D37CF22B3EB29400C45E5000C161250A040225662BF02FE98D6",
            INIT_RAM_14 => X"2016DB528401BC1B31089935A880991602031CB2016C32040CDF193E8200488A",
            INIT_RAM_15 => X"C9BE7DDDCEC45069CCBE50C429BE506ECA3FAA156040A204D942536D920008DD",
            INIT_RAM_16 => X"962428A4C940CFFAC08EA2852A2A25AB0C80525581438E71F62A61D3BF72059B",
            INIT_RAM_17 => X"4A40195556EFFC488C732D5A852224C889B340095CBC508A4199066D714D34A8",
            INIT_RAM_18 => X"8CC93C708006AC721B862318602C01212258D2CE44080C0911B7FFE488384011",
            INIT_RAM_19 => X"1664B20582486B096DC93F761554AC21ED5A1832824B345B423A3401565022D3",
            INIT_RAM_1A => X"E39A83371278E663BC0B1BF1E5E1000D2436C540240078096C03664B205992C8",
            INIT_RAM_1B => X"25311085A8A28353CC9EC427B10012FCB7ECF51905B4349160D5C48CB20EA029",
            INIT_RAM_1C => X"422B02856A0C0AD1CA3495D96324C224420C4208C200C2A15962E86D50CD21FC",
            INIT_RAM_1D => X"F056013D840BAFC5BD89015A00028449C55865048F8D12B483CCB84C224D8C69",
            INIT_RAM_1E => X"5AD625192CA1B0B2EF37EA310192F34A325946F20F4CD1DBB456EE63C1999820",
            INIT_RAM_1F => X"52D00000019FE208805BFE601398005F7A9801BFFFFBFF730FFE51772412ED29",
            INIT_RAM_20 => X"97B6A1C61A005A50A952155B13C5545DD3BEC93BE9D969D8A0ECD699493B0999",
            INIT_RAM_21 => X"3662D18D53B5529C6B462D904030410F2987F76AE99082301A76DFFCDBD280F8",
            INIT_RAM_22 => X"B9C0D70012C8100F02A57E94F585103548FF1A788E13666C0FB4D30C24833694",
            INIT_RAM_23 => X"A5449038F03B7FEE480307F1102CC52451C0C25B0829B0EEFDE03D3D04142A51",
            INIT_RAM_24 => X"1854A05040027D0002B7F59B59C74C1766AA3151C10A1F5823656671E023EDE4",
            INIT_RAM_25 => X"F1D0AF734000640F8BAD82B5BAA3880AC05C0BDC7B96FE9AF64C00BA23C80332",
            INIT_RAM_26 => X"8324E2621D8F4B2578AEE658FF1EA65185D11F0800600588B1001801688C402E",
            INIT_RAM_27 => X"DA0F9D292022728848197B2E8F96145887303588887D43171EA08207E2C32C08",
            INIT_RAM_28 => X"A3D5A2576AABAEBBA1EA5AE10DAAD52414511401400DADA8096002B29A3DD539",
            INIT_RAM_29 => X"3726B597AA78A800C841394877FBFFFFFFEFFFEA95559D4C16AFD65F97EA7A28",
            INIT_RAM_2A => X"6A1347C1D90061090065BFF375FDD0F8E988E4274031B1887FC3E66678809F45",
            INIT_RAM_2B => X"000F6677ACE21AC02FE7209AEDA8CB4201B4F1766126054967611195182E7D90",
            INIT_RAM_2C => X"8D662F3EC87ED1491AF32277F3C0BB100148622E0CDF73EACE41E12A61721B80",
            INIT_RAM_2D => X"A99736C201F09D0F807491FC11C7647DDB62BB24B293E68999B65D7081DF3252",
            INIT_RAM_2E => X"808272F5F5A954A45BB83A775740002AC682D4010C5355C23772E82D0FA87E35",
            INIT_RAM_2F => X"29AE35540024894036BD6D5B6A48126C0254A5FC845007121155575652C0B774",
            INIT_RAM_30 => X"62280010246122210C8D050D801929C3A10032DADD79E0AD0A48282D89E28C59",
            INIT_RAM_31 => X"10A8A09916C82645B26C932582440590706C92449B24912012A008075E01882C",
            INIT_RAM_32 => X"F1F78129454A607B0294BDE97ED3640C5746110020B09020826699949A044181",
            INIT_RAM_33 => X"474C99DFB9715D37CF22B3EB29400C45E5000C161250A040225662BF02FE98D6",
            INIT_RAM_34 => X"2016DB528401BC1B31089935A880991602031CB2016C32040CDF193E8200488A",
            INIT_RAM_35 => X"C9BE7DDDCEC45069CCBE50C429BE506ECA3FAA156040A204D942536D920008DD",
            INIT_RAM_36 => X"962428A4C940CFFAC08EA2852A2A25AB0C80525581438E71F62A61D3BF72059B",
            INIT_RAM_37 => X"4A40195556EFFC488C732D5A852224C889B340095CBC508A4199066D714D34A8",
            INIT_RAM_38 => X"8CC93C708006AC721B862318602C01212258D2CE44080C0911B7FFE488384011",
            INIT_RAM_39 => X"1664B20582486B096DC93F761554AC21ED5A1832824B345B423A3401565022D3",
            INIT_RAM_3A => X"E39A83371278E663BC0B1BF1E5E1000D2436C540240078096C03664B205992C8",
            INIT_RAM_3B => X"25311085A8A28353CC9EC427B10012FCB7ECF51905B4349160D5C48CB20EA029",
            INIT_RAM_3C => X"422B02856A0C0AD1CA3495D96324C224420C4208C200C2A15962E86D50CD21FC",
            INIT_RAM_3D => X"F056013D840BAFC5BD89015A00028449C55865048F8D12B483CCB84C224D8C69",
            INIT_RAM_3E => X"5AD625192CA1B0B2EF37EA310192F34A325946F20F4CD1DBB456EE63C1999820",
            INIT_RAM_3F => X"52D00000019FE208805BFE601398005F7A9801BFFFFBFF730FFE51772412ED29"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"073FB6073F0040B92E0CBD6351C97B7A096D85D65A9A70A08017FD0101010715",
            INIT_RAM_01 => X"6D35BBC80D7AAB45F7D6925B0C85F631C1F584CDD01D702873D8A5FAE92FBBCF",
            INIT_RAM_02 => X"9C40F6273B91F19228FBB1C30E529DBE24AAF381965DD401755420A42BDCB296",
            INIT_RAM_03 => X"2170BF5703010918DF57E4D5C8705655F23773EAC3900E2074BD5BAC7C2446A3",
            INIT_RAM_04 => X"A0320D41106A01033646F0C02FF8C145100143D24CC6A6F8838A404CC52D3088",
            INIT_RAM_05 => X"12F2E641F7D594B6F29781050E94203AE0CA8D4330119AC5AC4759488C18420C",
            INIT_RAM_06 => X"FAEBF94EDC42442419779CB2FC00A0F1356A65F2DE00A513047343ABCC802082",
            INIT_RAM_07 => X"7CE9EEE63315696CA351BA4406555C822088246AC51A351BA440624104026743",
            INIT_RAM_08 => X"021E6C1106373CFB57911FD4C9EFAEB6DCDD76BB099832A101EB7A7E5BA8D64F",
            INIT_RAM_09 => X"0AA00A00296DA4DCCC4554C4A024013E969DE223A1188F28807374038B84A5E4",
            INIT_RAM_0A => X"AE48B924364488CC29126B8D3218A9AEC135838B210041F7C04244F8E09215C2",
            INIT_RAM_0B => X"2DD6ACE743B72B59DE43758CFFD409813C94381C6698049E4562631B010AFF74",
            INIT_RAM_0C => X"62890BBC88470A0F50BDC8DCBA89FD4085EB3A2100B005DDEBD06839937A86EF",
            INIT_RAM_0D => X"9432C451407EA5E39001024863D080285F23DA4007721690F082F8E25F7D2280",
            INIT_RAM_0E => X"1D904D809267D8218A1AED111678101084A5508F79D84A784FFD77AD720122A2",
            INIT_RAM_0F => X"EB8DCBDE72033EDAC8C5151FD76CBC450B2CA516DE9331DA383A3A3A383A9211",
            INIT_RAM_10 => X"011400003FEBBF8541BFD47E4ECCA516DED76C2EAB6504259FE72029280008E9",
            INIT_RAM_11 => X"3C7AF06624218719D00CE1C9292545FE924A8054050504114411415541114144",
            INIT_RAM_12 => X"500BE7C2F1B14DCCEDB16083B81FFDF02E5F42D2F85A3EBBD6B975AAB1FEEFDE",
            INIT_RAM_13 => X"5104975A3707A41440306F8A40494A24EBF3F33D1D6ED7C65BCDF5AFDD27FE2D",
            INIT_RAM_14 => X"25050F66606510512871D91B9D90EE6C80530DCD988E82CAF72A802D407B9998",
            INIT_RAM_15 => X"87333026740483349B221B72020E11F9807512086A12CF33707E28937F126256",
            INIT_RAM_16 => X"BEC5402B80E87B80397A20450C01012C848C91400112484603E5599731048811",
            INIT_RAM_17 => X"329732E76C2DAD8F19DD7D4CB675B39FB47D29BB7B0A6F172649434CB5FB00A6",
            INIT_RAM_18 => X"C6B19C3CC2CF30B6D9CEF3151354E666F975A95223D0B8CA4E167804B4920687",
            INIT_RAM_19 => X"5217504E59BB980D9B7A84CDB6D200A3592C4A526653FE37F058391BA860CE20",
            INIT_RAM_1A => X"1B340D4679C99FABCEC8C7438D3CA8198BDC28E20B204583014908B32C60B51D",
            INIT_RAM_1B => X"6AB82D2A0A1D440AF72D421CC444C84D8B77D540A81DA85A8130B64D06CC22D5",
            INIT_RAM_1C => X"6F53A00ECB92CB70B0F2E4100107E33424A6EA05056F5283841A941DA8669505",
            INIT_RAM_1D => X"241810039410003412280290992D03BAAADB25EE7041C965A0511C90F40601E8",
            INIT_RAM_1E => X"698A010C960500681E9100801A003241800E50100201A291400068100A41A183",
            INIT_RAM_1F => X"94251D3456C3CD102D898003BAAAD85B1385B2811DAAAD45205AAD6A3580C0A0",
            INIT_RAM_20 => X"08402F450805C39A014E17830065724A432AB6107B7D920840D10920D1208674",
            INIT_RAM_21 => X"8E354086846A1CC4D438CC882CEA10E6C7B02AA4A427CAA1161FF80000A81042",
            INIT_RAM_22 => X"BB4CCDCB2CCCCA2BA603CB67272644C45D8823DAD4EE264643941853F354CA7A",
            INIT_RAM_23 => X"A48A9B32B19A00E2BBAA5E898408A6E52007DA5161520115CB8881590A96E584",
            INIT_RAM_24 => X"7347537EEDE66FE65C88D8E4E3360E18405111646C8686EEEEEEF18AB2226341",
            INIT_RAM_25 => X"06CB3C1A97970787E16797973020EC2DEF5C128D3F93266DAD483A1F4F598908",
            INIT_RAM_26 => X"00514CB58616252603AC378859B63030632931442D30498B052B848AB3032F21",
            INIT_RAM_27 => X"06A608309B8C68153D2D4AE30C8C480A8C26A5102055C806DAA25E31FC32BC02",
            INIT_RAM_28 => X"7BF1F0F80102769DAD77B20110D0BF048F8183122461707F8D84E6D588ACA4DA",
            INIT_RAM_29 => X"64BBE0004F075B296E605BAD94AE005B38CE804647091002E7C3C170C327A100",
            INIT_RAM_2A => X"D05BC303381E587AD105183D6C82601300A3062D999C1CB28A64470441ACFF53",
            INIT_RAM_2B => X"D61D60E018032220437C820979C0180C4D336B1CEA3102C8591048C189108130",
            INIT_RAM_2C => X"FFE83B25EC064D0598DEFA829180DC0399C0391B09600221AC00759D4A0EA041",
            INIT_RAM_2D => X"303364B2B14C18D83039C5A68CDB2066D4C61BE1DD87731110A2C28CC418AD85",
            INIT_RAM_2E => X"00000C022382049003603FF0916500708A153588CACB8963C4C31C6C0292CA2A",
            INIT_RAM_2F => X"E044C9D3012630D00A83C00196F310703C4804A3704EE088208010C838000000",
            INIT_RAM_30 => X"307678687820040814254582B009C18185C2C64B241AC60006174982B00184D1",
            INIT_RAM_31 => X"488C448A253DC0E0EA0140BF613E44443C8A089508C43A898ECCF07004A21130",
            INIT_RAM_32 => X"0A84B1550736DBF40D0594532F3CF22C6F07007E2C8D6387679647594613C040",
            INIT_RAM_33 => X"A3949DFA7FA36C909CC2244C192211991390142C2800094242C8880089CC1A33",
            INIT_RAM_34 => X"18064172563F53228E9324A52828DF04A86184019204E0404A3A49A5608E7AF0",
            INIT_RAM_35 => X"22B1449D69D5A25D036E797B0296B204D30201B48BCBF3C2379167CDE0800900",
            INIT_RAM_36 => X"37F418AFB3D591B2668D8C329723839A376C5A7941A002400C1C00C1C00C1C04",
            INIT_RAM_37 => X"4290709ED40840DB9B1C6B1083402104806170CA64041083497ABA0280D88913",
            INIT_RAM_38 => X"229FEA8F0C70D7D217EFE59B1679E4FAF618686B0258C406C9C30442004807FA",
            INIT_RAM_39 => X"57EAF7406B851A2C0A582C252ADA624651FB98731D9B7351A80B7739A896E0BD",
            INIT_RAM_3A => X"480214E09F22BEA53A49E7B24EDFC6A021100D4154DEA72404E0AA5E41D79F67",
            INIT_RAM_3B => X"0740F407944CC4998808FFFA519600CB4C0E9E93298C2265B793DE07150500EF",
            INIT_RAM_3C => X"92118419608A0630B0109832C325961054CC86CBA2CA9F5594A2AD1CE6666660",
            INIT_RAM_3D => X"88E8824D1CB90ADB735899370C828961811F9106111930C4463CC45827303431",
            INIT_RAM_3E => X"DB4ADA5EC9A7DCC78E8FB8C736994B60F9B8B71934884462268AA504D49A75FC",
            INIT_RAM_3F => X"169A1B623A7F15AAFDE4E46C6CE4C804ABD4584D3134C05F3C9D4D8ACAA982ED"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_2,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"AD5751BD429B4F61318427560CE39D492990013FD212081064E2FFF009FB997B",
            INIT_RAM_01 => X"8C6AC955A8A6140421573E413CF5A80AA1436D8B4C31A2AB26D2A61CE834248B",
            INIT_RAM_02 => X"6CDEE7468681D6C31E4991CA3736E9ACB7531EC6D8BBCD453718101EA25D7927",
            INIT_RAM_03 => X"15408676F600F490FAA59B488C7998CC8CCC28922AC62644EEBB432EEECB51B1",
            INIT_RAM_04 => X"DDBB7B207EFA17098E07684801BD45625A36BB62220506E171891964A31BED22",
            INIT_RAM_05 => X"FA4F91915C6AC9D8570C292F10848189906127BCBE06FFE92DAFB4AAFB240D88",
            INIT_RAM_06 => X"4CA272352720BCD900A6D79BFD9D0595EC0D044ABC8CC28E9AE946E3D2000A4E",
            INIT_RAM_07 => X"9C8CA06AA05B63C89A59A3E4E80807B27A70B0006624C4AC4A0995CCD8CA2082",
            INIT_RAM_08 => X"06C78011F78D8B82E59F0CD4B32D6801669BE3EB0B96960DFF152005EC7C16CB",
            INIT_RAM_09 => X"3AE624C94932927924D20024CD638A01C8620023319662D80E05805625BC4A40",
            INIT_RAM_0A => X"8366123AA809AB30B47977571C5D70397A93C723106D0A2C254714359DC7C9E1",
            INIT_RAM_0B => X"39BCEF6BF4D23532957455F1C80115524179D59C4C5D34DF7296991146CE2450",
            INIT_RAM_0C => X"9E2DBCBF62498A769883D7218899245CD18AE49F0146517422EE475D520029ED",
            INIT_RAM_0D => X"E9969472A81B83113144528F831AA6C3221E137C1E9C670E26808A894013828D",
            INIT_RAM_0E => X"9FE2D1F27443253D58403577C801AE23371F00290A17E1C4A40258BFD204230E",
            INIT_RAM_0F => X"20721F982534A8179F13E2C6328CDE7D2A73087D3A9314419022103DFF767776",
            INIT_RAM_10 => X"7DE6C2ED45D76325CA2A8E198859334553AB02945CAB1F17C142288008073004",
            INIT_RAM_11 => X"0644C9567C0BF9911B870B989C59330089AA4C8065AB1B11132213EE0FD83081",
            INIT_RAM_12 => X"6AA394A8644494895569192AE42AB508290A2CA59B4D6EF213548EED8642F231",
            INIT_RAM_13 => X"71163594CEC5863F0F56625E221D6B8180848C6B2BE24CA2AEEE5D187201CAAE",
            INIT_RAM_14 => X"198817644F293AC1946061117122A39D8841818C1389D51BDAC5491819025165",
            INIT_RAM_15 => X"27929938B8E10530250877A4998D0DF0004852125C20CA8D4279881E41208B14",
            INIT_RAM_16 => X"5E1384C93920A16C9B696272DE7A2948BE8AFE81310146B8AAE5E549FA27EFBE",
            INIT_RAM_17 => X"376E511217E00B624A46BA2E4CC10B729C326F710F24CFE78C5E63F3034737CC",
            INIT_RAM_18 => X"EFD5995634050D4CFEC166B032BEED5553AF0358304080D9DD0A2E9948593830",
            INIT_RAM_19 => X"C80CEC08A7F5F85CE65326632B4C4F3920019A35AE2AEB3A1131046EE45B81D4",
            INIT_RAM_1A => X"5939FC47C933E1B0AEF12AC84454CA47B00A6BEC5402AA08B5106E3065602454",
            INIT_RAM_1B => X"EF40312A73337CBAD4838F42A32938588D169240D8E652F6D72D8D19D56DD767",
            INIT_RAM_1C => X"E2E0440C6CBD60741FC178643A852D4A2A0627C688D905B882524E191E7951EA",
            INIT_RAM_1D => X"36E0548D65FF9125A765F0220F6EB9D1B318244CC6CA2CBC9CEC6979C14EB28D",
            INIT_RAM_1E => X"082C891C76A4845096304A0D8502080C1198921998821D11C29CA830C3374992",
            INIT_RAM_1F => X"35C65240B61076066A23CE4CFC5E76063A1C2AE07DF555007338BDC080EA0C23",
            INIT_RAM_20 => X"639303AE5376F664C7125632C19440CECD5740C77849D937472B202579964F60",
            INIT_RAM_21 => X"14E5DCCAFE50CC13922A5B149C598A621F80C24D215291228844E7F33F9763C6",
            INIT_RAM_22 => X"21D9DC46629BB376E97F2C7BF8C3A218EE79DDBCF886B2BBDE702F71B38AEC69",
            INIT_RAM_23 => X"6EE48A1CA6430860DE613153615CAF4C8D191004CE9C6105D8C6795B6484467D",
            INIT_RAM_24 => X"9F0120108829220B230F44550832C1022530CC13C4C30D8254ECA5200A194126",
            INIT_RAM_25 => X"C0BED5FBD379F904A41BAFB6BE4EE9F6E8058229DD0C354F03CA6C4D8B6C16A2",
            INIT_RAM_26 => X"5621E625522D34519BF2C353F8AA030B9109C2F9686AD36F57AF3016D9160354",
            INIT_RAM_27 => X"5FFE6AD3343986C4103935236B6E6E11B940EF46A8FC06E6872A6929D50DCDB7",
            INIT_RAM_28 => X"7740114D6B08228BCC693FB12CECCCD2461586069445ACFC910B1241434622B6",
            INIT_RAM_29 => X"C08C4847914664518E27EF7EB9C870A226AFC35BEDB651840466400D4B3C0F87",
            INIT_RAM_2A => X"A807C3A1110211AFCA2A142F0BA928156D142250438143D339E4E2079F298493",
            INIT_RAM_2B => X"7FF29C990C9E66273CC78041192D03081CC62A8A0D8CB4D9CF2F2558131A78B8",
            INIT_RAM_2C => X"527CCD419525AD29AB7D372C0B56AA0A065F8BDC905346478059EC8280192068",
            INIT_RAM_2D => X"12D552A8A0496EFE3AAC6F34739A94E798101823148D811212E9A349CB219049",
            INIT_RAM_2E => X"01DEC1A54696B9912E8B0705C8587D4F7D36C863897BD3102AA663B819B55B7A",
            INIT_RAM_2F => X"2C05EF54A3C0F7F5F017E03F5800377CCF6E493C84E8F56441831087370A0848",
            INIT_RAM_30 => X"100E0A7211342DF02958046899EEBE6E491299A09312778193FF3D7FFABA8000",
            INIT_RAM_31 => X"1A94A248414CE030020F207BF040A06A3DF993DEA3823423F405294A52014565",
            INIT_RAM_32 => X"AA0AAA22B1C70003F542A66FD1F1CF9D4578315F8C1C6FEC4FEDBDF22CB20482",
            INIT_RAM_33 => X"00D988737BBB44C414210118C673B0C1BDF76C499226F78FF41A0AF7AFD3308A",
            INIT_RAM_34 => X"6087F8B130F04418C0A1C082FC005843F5B42CADD9455ADBD328C13219110DE1",
            INIT_RAM_35 => X"54E09A38775020189010680840800297C31282442326D008D1F2351A89FFD7C1",
            INIT_RAM_36 => X"A0D8E36A84D5C61285128845215F8F8821C308E368283D8E2B42989C04A8B513",
            INIT_RAM_37 => X"81F3167814687CBD683E54D44555E6C95B5F2A72C0C193C6110C0221A448D0C9",
            INIT_RAM_38 => X"C81822450A1241244495470389D430FE8DAA04503442C4F91309238ECB252072",
            INIT_RAM_39 => X"C2CAF43524E5545491F070E856F5E4B404415ED956AD5A2A6A6B0016961D4697",
            INIT_RAM_3A => X"AB9930C7AF100009166F6FB3DA3EF3FB9D1A2C03ADCC009791FFE793B301F7FD",
            INIT_RAM_3B => X"8000000040A7AACEB6957E89D7F588DAFA30E0194271568A533159838C696997",
            INIT_RAM_3C => X"000000000000000000000000004891883F511C904DC134F4DFC5FE73F7DF2493",
            INIT_RAM_3D => X"0400280000003C3406303220344C403C04001000101000000050627424000000",
            INIT_RAM_3E => X"80000000424202423E1E3E02304C3C0C3C7E7E40403E427E3402421824347C1C",
            INIT_RAM_3F => X"4200000042000000000000000000800000000000000000000000000000300044"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_8: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"10B2E5DF7980090C232ED509694969961C60E62090182066C2E6CD3676DAB088",
            INIT_RAM_01 => X"CD2B852F6B6510104A08A2ED5469061B9B28C9CE99D8E8F006F6D46C62FB8011",
            INIT_RAM_02 => X"2BC21E09C7C864019BB96E98A1879949C0DC07BCEF70B3930C9B31F30CB1D9DE",
            INIT_RAM_03 => X"255CF189100C982AD03DEBFD9F92C5B459C37BD9B9ADB8FA0C130C8CAD016144",
            INIT_RAM_04 => X"18BDA9E802F38F0002BCFF9151C74C2B72BA01CC165AD1585B38890DC25D59FF",
            INIT_RAM_05 => X"F035BC14D410AFAEFFE82CA5362D086485EB4C185BDED4C387062C24B763E777",
            INIT_RAM_06 => X"8B78E66B68B4899002A44440557D96FE2125BBE3E445C052DC79117012D71E20",
            INIT_RAM_07 => X"170ED531F23A03CA7911723ECD159708792E7DC1F35B42F702F18A96AEB0EF08",
            INIT_RAM_08 => X"998C02352E7451426613C2E30887D586987194099FC5828124EABC32A665CAA8",
            INIT_RAM_09 => X"6865975639ECEB973D7CCCEF9800000000100016C000694580405CA1289A7A1B",
            INIT_RAM_0A => X"4F173EA5F0E710FFF9159993FFF7D66CBEE261883F4E6E837973B9D9903491E5",
            INIT_RAM_0B => X"10A098DFAEBC9ED53F88479AC32E7E6D2E39D9DB4E99E2EE5C3FBADD9720147E",
            INIT_RAM_0C => X"8E29939936952D695C49987F8014128AE912C7C26664CFDBB3F135D98174C8C0",
            INIT_RAM_0D => X"FDD50657043241919F04423A8F0491BD8973C3C311CCD8C9D8CDA4C6DCD989B3",
            INIT_RAM_0E => X"95BFA2FCDB7FF24950EC1A3D9F87022E9783EA99EC62FFD2EAA82A1EA0EFDBF4",
            INIT_RAM_0F => X"9DBF3FF87021C1E6ED028BAD9B697F936BAE900A49755F610EAAABD1A576DFF8",
            INIT_RAM_10 => X"99CE19CF147D3D31876585EB49213DFFAC93B8C89909A60F70EE403D9582C051",
            INIT_RAM_11 => X"1298F524BB6C6DA7FF7ED9B7CD07C3FC7736D8925FFEB6D063B8E789660667B0",
            INIT_RAM_12 => X"E0B88519E12A994CB7BDE73000B9BE207A14C8C1265CC84439DCD1E4F132C101",
            INIT_RAM_13 => X"8760DD83197B9D368E4AC4003E80F33786C824CB99519C6DC9C763C1080484D4",
            INIT_RAM_14 => X"324F7FEB6F05B73B1DC39DDAE54A64D31603DE3ACF283C3C22C9EFCA86A642D2",
            INIT_RAM_15 => X"E03070596F3A687D6C2BE5A1E6678990EDBDFA35FC5CF793B9D96DFFFBF9F417",
            INIT_RAM_16 => X"5980B2C20D96B00064A263E499BACFFE10A07BFF0DF7A76119CD69F9E67C2D24",
            INIT_RAM_17 => X"4C31D1F7FE9D45192B52F72E732B36E4AFDB230FD4D7196C5B1611433BE47E39",
            INIT_RAM_18 => X"0B2A7C49012FD3FA5D891B997108CBF7D96E437856458E5FFD075574386CC161",
            INIT_RAM_19 => X"6936F89343270467F37CC634D34EBE0E0489081E7836A092418108C35FC83ACA",
            INIT_RAM_1A => X"787666B8DB9E1D611CAF6FAF1EDD001E7F3FE74009EF7CDFB6B4936F8935FF6B",
            INIT_RAM_1B => X"05B4129128A20208D3A8F32A3CCAB8D67745E9DAF5E6C67A582E36EAEB11A0A6",
            INIT_RAM_1C => X"F7AB8BE36B8D88B106A011C4A304C32C43284600D602D2837502EC7450EC61BC",
            INIT_RAM_1D => X"FC17812F0F0B436D55D501BB42C4270C0578915C883BAAD4E1B158AC55B25A69",
            INIT_RAM_1E => X"5EE776E7BEB63D3EFFC1B5BC29383BEDCF7D658A8C0CDEC334D00004A7FFFF70",
            INIT_RAM_1F => X"70000000027C79AA91983EC0DF180500008A0CB5810B56F3BAF058041BC68054",
            INIT_RAM_20 => X"10B2E5DF7980090C232ED509694969961C60E62090182066C2E6CD3676DAB088",
            INIT_RAM_21 => X"CD2B852F6B6510104A08A2ED5469061B9B28C9CE99D8E8F006F6D46C62FB8011",
            INIT_RAM_22 => X"2BC21E09C7C864019BB96E98A1879949C0DC07BCEF70B3930C9B31F30CB1D9DE",
            INIT_RAM_23 => X"255CF189100C982AD03DEBFD9F92C5B459C37BD9B9ADB8FA0C130C8CAD016144",
            INIT_RAM_24 => X"18BDA9E802F38F0002BCFF9151C74C2B72BA01CC165AD1585B38890DC25D59FF",
            INIT_RAM_25 => X"F035BC14D410AFAEFFE82CA5362D086485EB4C185BDED4C387062C24B763E777",
            INIT_RAM_26 => X"8B78E66B68B4899002A44440557D96FE2125BBE3E445C052DC79117012D71E20",
            INIT_RAM_27 => X"170ED531F23A03CA7911723ECD159708792E7DC1F35B42F702F18A96AEB0EF08",
            INIT_RAM_28 => X"998C02352E7451426613C2E30887D586987194099FC5828124EABC32A665CAA8",
            INIT_RAM_29 => X"6865975639ECEB973D7CCCEF9800000000100016C000694580405CA1289A7A1B",
            INIT_RAM_2A => X"4F173EA5F0E710FFF9159993FFF7D66CBEE261883F4E6E837973B9D9903491E5",
            INIT_RAM_2B => X"10A098DFAEBC9ED53F88479AC32E7E6D2E39D9DB4E99E2EE5C3FBADD9720147E",
            INIT_RAM_2C => X"8E29939936952D695C49987F8014128AE912C7C26664CFDBB3F135D98174C8C0",
            INIT_RAM_2D => X"FDD50657043241919F04423A8F0491BD8973C3C311CCD8C9D8CDA4C6DCD989B3",
            INIT_RAM_2E => X"95BFA2FCDB7FF24950EC1A3D9F87022E9783EA99EC62FFD2EAA82A1EA0EFDBF4",
            INIT_RAM_2F => X"9DBF3FF87021C1E6ED028BAD9B697F936BAE900A49755F610EAAABD1A576DFF8",
            INIT_RAM_30 => X"99CE19CF147D3D31876585EB49213DFFAC93B8C89909A60F70EE403D9582C051",
            INIT_RAM_31 => X"1298F524BB6C6DA7FF7ED9B7CD07C3FC7736D8925FFEB6D063B8E789660667B0",
            INIT_RAM_32 => X"E0B88519E12A994CB7BDE73000B9BE207A14C8C1265CC84439DCD1E4F132C101",
            INIT_RAM_33 => X"8760DD83197B9D368E4AC4003E80F33786C824CB99519C6DC9C763C1080484D4",
            INIT_RAM_34 => X"324F7FEB6F05B73B1DC39DDAE54A64D31603DE3ACF283C3C22C9EFCA86A642D2",
            INIT_RAM_35 => X"E03070596F3A687D6C2BE5A1E6678990EDBDFA35FC5CF793B9D96DFFFBF9F417",
            INIT_RAM_36 => X"5980B2C20D96B00064A263E499BACFFE10A07BFF0DF7A76119CD69F9E67C2D24",
            INIT_RAM_37 => X"4C31D1F7FE9D45192B52F72E732B36E4AFDB230FD4D7196C5B1611433BE47E39",
            INIT_RAM_38 => X"0B2A7C49012FD3FA5D891B997108CBF7D96E437856458E5FFD075574386CC161",
            INIT_RAM_39 => X"6936F89343270467F37CC634D34EBE0E0489081E7836A092418108C35FC83ACA",
            INIT_RAM_3A => X"787666B8DB9E1D611CAF6FAF1EDD001E7F3FE74009EF7CDFB6B4936F8935FF6B",
            INIT_RAM_3B => X"05B4129128A20208D3A8F32A3CCAB8D67745E9DAF5E6C67A582E36EAEB11A0A6",
            INIT_RAM_3C => X"F7AB8BE36B8D88B106A011C4A304C32C43284600D602D2837502EC7450EC61BC",
            INIT_RAM_3D => X"FC17812F0F0B436D55D501BB42C4270C0578915C883BAAD4E1B158AC55B25A69",
            INIT_RAM_3E => X"5EE776E7BEB63D3EFFC1B5BC29383BEDCF7D658A8C0CDEC334D00004A7FFFF70",
            INIT_RAM_3F => X"70000000027C79AA91983EC0DF180500008A0CB5810B56F3BAF058041BC68054"
        )
        port map (
            DO => prom_inst_8_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_9: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"10B2E5DF7980090C232ED509694969961C60E62090182066C2E6CD3676DAB088",
            INIT_RAM_01 => X"CD2B852F6B6510104A08A2ED5469061B9B28C9CE99D8E8F006F6D46C62FB8011",
            INIT_RAM_02 => X"2BC21E09C7C864019BB96E98A1879949C0DC07BCEF70B3930C9B31F30CB1D9DE",
            INIT_RAM_03 => X"255CF189100C982AD03DEBFD9F92C5B459C37BD9B9ADB8FA0C130C8CAD016144",
            INIT_RAM_04 => X"18BDA9E802F38F0002BCFF9151C74C2B72BA01CC165AD1585B38890DC25D59FF",
            INIT_RAM_05 => X"F035BC14D410AFAEFFE82CA5362D086485EB4C185BDED4C387062C24B763E777",
            INIT_RAM_06 => X"8B78E66B68B4899002A44440557D96FE2125BBE3E445C052DC79117012D71E20",
            INIT_RAM_07 => X"170ED531F23A03CA7911723ECD159708792E7DC1F35B42F702F18A96AEB0EF08",
            INIT_RAM_08 => X"998C02352E7451426613C2E30887D586987194099FC5828124EABC32A665CAA8",
            INIT_RAM_09 => X"6865975639ECEB973D7CCCEF9800000000100016C000694580405CA1289A7A1B",
            INIT_RAM_0A => X"4F173EA5F0E710FFF9159993FFF7D66CBEE261883F4E6E837973B9D9903491E5",
            INIT_RAM_0B => X"10A098DFAEBC9ED53F88479AC32E7E6D2E39D9DB4E99E2EE5C3FBADD9720147E",
            INIT_RAM_0C => X"8E29939936952D695C49987F8014128AE912C7C26664CFDBB3F135D98174C8C0",
            INIT_RAM_0D => X"FDD50657043241919F04423A8F0491BD8973C3C311CCD8C9D8CDA4C6DCD989B3",
            INIT_RAM_0E => X"95BFA2FCDB7FF24950EC1A3D9F87022E9783EA99EC62FFD2EAA82A1EA0EFDBF4",
            INIT_RAM_0F => X"9DBF3FF87021C1E6ED028BAD9B697F936BAE900A49755F610EAAABD1A576DFF8",
            INIT_RAM_10 => X"99CE19CF147D3D31876585EB49213DFFAC93B8C89909A60F70EE403D9582C051",
            INIT_RAM_11 => X"1298F524BB6C6DA7FF7ED9B7CD07C3FC7736D8925FFEB6D063B8E789660667B0",
            INIT_RAM_12 => X"E0B88519E12A994CB7BDE73000B9BE207A14C8C1265CC84439DCD1E4F132C101",
            INIT_RAM_13 => X"8760DD83197B9D368E4AC4003E80F33786C824CB99519C6DC9C763C1080484D4",
            INIT_RAM_14 => X"324F7FEB6F05B73B1DC39DDAE54A64D31603DE3ACF283C3C22C9EFCA86A642D2",
            INIT_RAM_15 => X"E03070596F3A687D6C2BE5A1E6678990EDBDFA35FC5CF793B9D96DFFFBF9F417",
            INIT_RAM_16 => X"5980B2C20D96B00064A263E499BACFFE10A07BFF0DF7A76119CD69F9E67C2D24",
            INIT_RAM_17 => X"4C31D1F7FE9D45192B52F72E732B36E4AFDB230FD4D7196C5B1611433BE47E39",
            INIT_RAM_18 => X"0B2A7C49012FD3FA5D891B997108CBF7D96E437856458E5FFD075574386CC161",
            INIT_RAM_19 => X"6936F89343270467F37CC634D34EBE0E0489081E7836A092418108C35FC83ACA",
            INIT_RAM_1A => X"787666B8DB9E1D611CAF6FAF1EDD001E7F3FE74009EF7CDFB6B4936F8935FF6B",
            INIT_RAM_1B => X"05B4129128A20208D3A8F32A3CCAB8D67745E9DAF5E6C67A582E36EAEB11A0A6",
            INIT_RAM_1C => X"F7AB8BE36B8D88B106A011C4A304C32C43284600D602D2837502EC7450EC61BC",
            INIT_RAM_1D => X"FC17812F0F0B436D55D501BB42C4270C0578915C883BAAD4E1B158AC55B25A69",
            INIT_RAM_1E => X"5EE776E7BEB63D3EFFC1B5BC29383BEDCF7D658A8C0CDEC334D00004A7FFFF70",
            INIT_RAM_1F => X"70000000027C79AA91983EC0DF180500008A0CB5810B56F3BAF058041BC68054",
            INIT_RAM_20 => X"10B2E5DF7980090C232ED509694969961C60E62090182066C2E6CD3676DAB088",
            INIT_RAM_21 => X"CD2B852F6B6510104A08A2ED5469061B9B28C9CE99D8E8F006F6D46C62FB8011",
            INIT_RAM_22 => X"2BC21E09C7C864019BB96E98A1879949C0DC07BCEF70B3930C9B31F30CB1D9DE",
            INIT_RAM_23 => X"255CF189100C982AD03DEBFD9F92C5B459C37BD9B9ADB8FA0C130C8CAD016144",
            INIT_RAM_24 => X"18BDA9E802F38F0002BCFF9151C74C2B72BA01CC165AD1585B38890DC25D59FF",
            INIT_RAM_25 => X"F035BC14D410AFAEFFE82CA5362D086485EB4C185BDED4C387062C24B763E777",
            INIT_RAM_26 => X"8B78E66B68B4899002A44440557D96FE2125BBE3E445C052DC79117012D71E20",
            INIT_RAM_27 => X"170ED531F23A03CA7911723ECD159708792E7DC1F35B42F702F18A96AEB0EF08",
            INIT_RAM_28 => X"998C02352E7451426613C2E30887D586987194099FC5828124EABC32A665CAA8",
            INIT_RAM_29 => X"6865975639ECEB973D7CCCEF9800000000100016C000694580405CA1289A7A1B",
            INIT_RAM_2A => X"4F173EA5F0E710FFF9159993FFF7D66CBEE261883F4E6E837973B9D9903491E5",
            INIT_RAM_2B => X"10A098DFAEBC9ED53F88479AC32E7E6D2E39D9DB4E99E2EE5C3FBADD9720147E",
            INIT_RAM_2C => X"8E29939936952D695C49987F8014128AE912C7C26664CFDBB3F135D98174C8C0",
            INIT_RAM_2D => X"FDD50657043241919F04423A8F0491BD8973C3C311CCD8C9D8CDA4C6DCD989B3",
            INIT_RAM_2E => X"95BFA2FCDB7FF24950EC1A3D9F87022E9783EA99EC62FFD2EAA82A1EA0EFDBF4",
            INIT_RAM_2F => X"9DBF3FF87021C1E6ED028BAD9B697F936BAE900A49755F610EAAABD1A576DFF8",
            INIT_RAM_30 => X"99CE19CF147D3D31876585EB49213DFFAC93B8C89909A60F70EE403D9582C051",
            INIT_RAM_31 => X"1298F524BB6C6DA7FF7ED9B7CD07C3FC7736D8925FFEB6D063B8E789660667B0",
            INIT_RAM_32 => X"E0B88519E12A994CB7BDE73000B9BE207A14C8C1265CC84439DCD1E4F132C101",
            INIT_RAM_33 => X"8760DD83197B9D368E4AC4003E80F33786C824CB99519C6DC9C763C1080484D4",
            INIT_RAM_34 => X"324F7FEB6F05B73B1DC39DDAE54A64D31603DE3ACF283C3C22C9EFCA86A642D2",
            INIT_RAM_35 => X"E03070596F3A687D6C2BE5A1E6678990EDBDFA35FC5CF793B9D96DFFFBF9F417",
            INIT_RAM_36 => X"5980B2C20D96B00064A263E499BACFFE10A07BFF0DF7A76119CD69F9E67C2D24",
            INIT_RAM_37 => X"4C31D1F7FE9D45192B52F72E732B36E4AFDB230FD4D7196C5B1611433BE47E39",
            INIT_RAM_38 => X"0B2A7C49012FD3FA5D891B997108CBF7D96E437856458E5FFD075574386CC161",
            INIT_RAM_39 => X"6936F89343270467F37CC634D34EBE0E0489081E7836A092418108C35FC83ACA",
            INIT_RAM_3A => X"787666B8DB9E1D611CAF6FAF1EDD001E7F3FE74009EF7CDFB6B4936F8935FF6B",
            INIT_RAM_3B => X"05B4129128A20208D3A8F32A3CCAB8D67745E9DAF5E6C67A582E36EAEB11A0A6",
            INIT_RAM_3C => X"F7AB8BE36B8D88B106A011C4A304C32C43284600D602D2837502EC7450EC61BC",
            INIT_RAM_3D => X"FC17812F0F0B436D55D501BB42C4270C0578915C883BAAD4E1B158AC55B25A69",
            INIT_RAM_3E => X"5EE776E7BEB63D3EFFC1B5BC29383BEDCF7D658A8C0CDEC334D00004A7FFFF70",
            INIT_RAM_3F => X"70000000027C79AA91983EC0DF180500008A0CB5810B56F3BAF058041BC68054"
        )
        port map (
            DO => prom_inst_9_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_10: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0E77E2373F00E88053194EB2101CB404828AD80900E4B8111126060101010400",
            INIT_RAM_01 => X"0B8646129B2413A20282672692421436DF494E662BF4B400E750204812000D86",
            INIT_RAM_02 => X"DB52D5BCF25BA0E824CF7770423082C0DA3B96BF478527E7A772A99F92E66CE9",
            INIT_RAM_03 => X"3CA0C94DA2D07393197D3B768BD35CD7E7634FDB84FC72F50F25309200DAC39D",
            INIT_RAM_04 => X"3AB45CEDD5644A9AC0574BA5AEA5BBAAAAEBF0011228F904A867884CCB94D664",
            INIT_RAM_05 => X"0ADD983DB6DF67675D29C101057342A3DC141442F695F8DF8DDF1CBEBD5B18AD",
            INIT_RAM_06 => X"7E7494ECD8204601D42D42672CF8121B2369A43C1DF234F20E0A903C5CF8674D",
            INIT_RAM_07 => X"70D10312604B5448CB65B298073A04B28B0A319A0BB8B45A298070514E42A957",
            INIT_RAM_08 => X"1B080C0616718F38C297BBF8AC02260B9CF49C4E0D9CAB090D1B09C6C024A8CE",
            INIT_RAM_09 => X"E98662CD96DA26FE667FF76CB6C7894022DF281EA0E830C08FF1222B0F062986",
            INIT_RAM_0A => X"E89911B63636EEACF816F16DAE8E96E96ECECE8DBECC01B6CDF77FDEEA0066E8",
            INIT_RAM_0B => X"FF3F2E97FBC7F15DEFE9CEC6B5138C60D506C7EA30080FF2254D231FE14B9C75",
            INIT_RAM_0C => X"2AC4CE326EF2CE8C4D796E97E26FF131AA8486C83D5D15719A4C29A4CFDFD3F7",
            INIT_RAM_0D => X"E0526AFFBF851800D070336C8C17FF3A71BC205E8002E26EEFB6071E8CE4EBFF",
            INIT_RAM_0E => X"191C7FF8FEC6FF48E96E97FFD7F8BA39D7BDBFF1A8DACA2CFF5D5E275244A2B3",
            INIT_RAM_0F => X"B843FD6A1A0D896EB674A335649C800B4FE697FC8BB2592DD5D7D7D7D5D4FC1B",
            INIT_RAM_10 => X"114144011500113BEBBBD501FFC697FC8B74BE23A5B7643720A1A0E9B741BEC8",
            INIT_RAM_11 => X"A54892EE21AA8B38D85573E8A5956355CB2AC001550054054105104451415541",
            INIT_RAM_12 => X"7C86005D099C4A270846BE4C47D2112F8608EA014908D7929F1F8EC34EB24E52",
            INIT_RAM_13 => X"01F7031B85653813DC512AB9113869EA060C91C81885782D264604F4228428E8",
            INIT_RAM_14 => X"876D363A723196DA69BB8EBDB8E8C3AEFC399874C18CE0D79D2439C12230E3A3",
            INIT_RAM_15 => X"10C0C3945A41A3AD342EF25988CB4CD10759FC6913D328C8C72B28DCA47D9DB9",
            INIT_RAM_16 => X"FCE74046C0A61BC2298A3051C2446204DF629452447383616AB9036C5820F333",
            INIT_RAM_17 => X"C2D17A666E046C7F274CB2F957736B1FB0016DA13291ED0C92D993F78DBABD48",
            INIT_RAM_18 => X"CE0240570BD5C2FAF3A23713E1CBB79856D5AE4BC3DB3B2536A827EE85D2A7D9",
            INIT_RAM_19 => X"7A7A489F9F6FE7DF3EDA4DF1249C42E705C9890111BCB476F9B17E7265DD56E3",
            INIT_RAM_1A => X"4B7C216B9B893CE91C38E737BCAE9FC674583AFDF4F3BA44FCF083569398A71D",
            INIT_RAM_1B => X"A1A92121FFE2B815F0F42679C64E484D29A2532A00B04C04C443496712D2895C",
            INIT_RAM_1C => X"4A2833FFFEFB6DCA1395F0BB7A822D380E452B30FFF1087FC0E843FE849090FC",
            INIT_RAM_1D => X"B7F123084C16020C4C90876DCDBFFD551F6DB7294FDF7DB6DEB399CB8AFDE090",
            INIT_RAM_1E => X"12C01FF648FA9C37FC200FB7F85BDB7F1C21300E09106064845C37F0F93FC03D",
            INIT_RAM_1F => X"D735ADABBB65EAE576DCDB55551F6DEDB87BFF7A8BC04002748040523ADB1F50",
            INIT_RAM_20 => X"C8BE18BEA07C082056E10C6DB788DB7DBC47DB3BF12FFD4FE0AEDB40AEA9A358",
            INIT_RAM_21 => X"7674BB9614266DCDCCD9D00927EA51FE9513E11CF03D411F427FF80030623985",
            INIT_RAM_22 => X"B0C2C8CB69D9DB3F460AAB2DC5B905B5576FAC671D6F9843DD2D644D01CDE9AE",
            INIT_RAM_23 => X"4CCE9BBEA52C295B4F08DED70036DBD3D00783200670E06E70917913BE9465CD",
            INIT_RAM_24 => X"3B5333786DC36F84580D8218F6D80D29755305C15650E3333333213ACE8A7353",
            INIT_RAM_25 => X"149EAB54B5E16CA55BB4D5E13F83303FE6F8D0E882892DB092A5291F4F5B3015",
            INIT_RAM_26 => X"0CB97A0E785D867D8BCB376AF017AC987BE36C579F533F0AD3FBB209CCB878B6",
            INIT_RAM_27 => X"5A320A5B49A94271C2F0026B6009369016D000DA60169216FF7A473F2B372B30",
            INIT_RAM_28 => X"D0BD309801A39E87F6CD2643C1B6EAD48D6362CC907228DD7963ABD762EB3104",
            INIT_RAM_29 => X"F98F385600B1EF9FCEE6F0F7CFEE86F0084F3EF5A7015BB0D12EB06BB0010967",
            INIT_RAM_2A => X"6E0F3058058886040760530203B01580EC1A6162286D910E58881B645D0C5741",
            INIT_RAM_2B => X"21931F57EAF21A0C5ED018C0554196E34F21E0C65B217A4AC15768F18B57B8DC",
            INIT_RAM_2C => X"11922EFF7B18F37EF0428B22C903581B6181B60F8340F1A0681F499258C90F19",
            INIT_RAM_2D => X"207372A2E36808DDA921D5A0CCDDEB84E18FDEB33545E6C68560B430280F7B6B",
            INIT_RAM_2E => X"00000C183F9AC69672D1E7E3593BCF5C8BA5358AD2CB696336A2D34B1392DA33",
            INIT_RAM_2F => X"B61CB9208F25CC23B8DB8078F10CD650306E459B5BD8B4AE4A9C6302305C0000",
            INIT_RAM_30 => X"5B414E7DCC2105C150E56672A0696761652E55CCE514340EC594897A8D8567DE",
            INIT_RAM_31 => X"F0BA57AAB23EB6A0B071FC6A5B2AD675286BCD4C694172DD0827AE70C435072D",
            INIT_RAM_32 => X"1A8FED4108C02409C90120B7A8431E889AE70C021A10B03818F71C0906BB8039",
            INIT_RAM_33 => X"A7C1D91A46367A6514D306481122911917C2B2983C141D4016DE8BBDA2CE5D63",
            INIT_RAM_34 => X"604D052256149DD7BB4A3485B6AEB016B7EFBEF14CFFB5E11EED1DB066C870ED",
            INIT_RAM_35 => X"A2C2449A5DA5F65248B37EBF2D46E80D9EF8D0EF9E7003D9EDC04D8D6E2ABD15",
            INIT_RAM_36 => X"3804362FA2DF5561D5D56B12E7334954A42B7C8C406781CF0696F0696F0696F5",
            INIT_RAM_37 => X"4212F02E96A85CBC7EDBE6810179021696715FCDE050C11B496ABA80FEBB0A15",
            INIT_RAM_38 => X"E00A014AF00C3823B710060708501D5E2BD65D2A0F18940CA30E401E12400FF2",
            INIT_RAM_39 => X"08005894B320914F0E5600D8E0315B3829451A632B315B8C045A6751A2903C23",
            INIT_RAM_3A => X"730BD4B915CC3A61BCCDF7E66FDB3216A11101B544C8CE7190C02134620D6280",
            INIT_RAM_3B => X"2440CE11C939BA737708000B59949A7169A6DB384FA9C065355D15B841C91029",
            INIT_RAM_3C => X"E299C7E670A2FDEA35B0CFCD8491F6ED9B1B088B4A8A4255C6A5509804E4E4E0",
            INIT_RAM_3D => X"56956C0DFE6ECA59364C9BA7F368DCC1E612854C2A26EDB227F80AB74CD591E1",
            INIT_RAM_3E => X"32B395BCAD5B0A5B35329485D6A68C7A3C1A7531F8DA7F773623B1ECC65B94F5",
            INIT_RAM_3F => X"24011A703855D4A815CE4ECEC6CED765C4480193C2DCF8C0B6B95367B6476333"
        )
        port map (
            DO => prom_inst_10_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_2,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_11: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"9E28CC30C7C2553DED3378D655AD194B2E6C1CFFED700F6713D9F8F33EFC361A",
            INIT_RAM_01 => X"71A553CCDD8ABA79BD27B7AF735ED2D34F1EF3A81A160C9ECB1B1FAE6EDEEFF9",
            INIT_RAM_02 => X"F6369572C3BB8AA1984A8D12F776E224ECEEB21F97FCD6C0CF17A044EC2BBF05",
            INIT_RAM_03 => X"E51D405CAF70F622DD4599602D7910DCAC8214B2A4202510C593202C8B164C8D",
            INIT_RAM_04 => X"34ABEB9DFAA4853910C9965C158947081CA41402E8E65478737F73BB629AAE2E",
            INIT_RAM_05 => X"F84DBBB9878C55457324E92D3DAE91D729AC76BBAD4C6EECA74DAB5EE9A175EE",
            INIT_RAM_06 => X"D7779D7B79D1C75DF87378E98719C1AF38B1B801C71D180CE86370AE9C2BF38C",
            INIT_RAM_07 => X"973FED2E9BEDBA474B70B121A8D60F3B4EE3F1A238FB3B730EDAEE74EC632DB4",
            INIT_RAM_08 => X"27271C28420E47B8DEC74738FC3EDF9FBD40EC09FC7B4D3A1475BE433705FB5F",
            INIT_RAM_09 => X"3091900604017933442359491FBAB63F346F0C5EC8E3A531984B09E605A30A06",
            INIT_RAM_0A => X"5699692496359B8E67A7E74D9A0FC504C8465638CF74A1AF9185921A7D262989",
            INIT_RAM_0B => X"352CD1DAFC910CC504334DF9E6F1F4F30161A36293C85CCF1CA13994ED29D34A",
            INIT_RAM_0C => X"F00030AFDB7F22E68CBAA4D9BE7633D3B53E90E4B124422A2A4454BACA5A8DC9",
            INIT_RAM_0D => X"D195D748900C29DF7F381280A9738CDC3BF5BBF937D3A4D99CE2ACCD97CEF2C7",
            INIT_RAM_0E => X"F1A8CCFC0C7A15BD9E7C2557CB00BF2584E16AAD13D7EDB525A85ABF90C0136D",
            INIT_RAM_0F => X"386BA04EF97A3F8551DAD9D24A8D259A03ECFF5AB81B1C31DFDAE10100544F8C",
            INIT_RAM_10 => X"7D94E6ED80D6722F3989B91E31C63B64C363DCE71A861C14382E270FC02878C7",
            INIT_RAM_11 => X"293A130C900FBA4EA70D2BA25B343C5B026D8E8766A4E4267CDAEC99E830D230",
            INIT_RAM_12 => X"3B9DDFE4F83A56E124BF5BCE9B34FCAA67E49B3A42E19184B6C9F07349210436",
            INIT_RAM_13 => X"B755D1CBF0DCF6FD40BEEC16EAB4A6D16839C98CBE9DA342FC69FB709F8E7999",
            INIT_RAM_14 => X"5ADFAF6726384795A7656B753D2369B9EB5595BAA722012DF8DCFBF15BF46D6E",
            INIT_RAM_15 => X"3AC884B1E69101135CD080022451F20884CCB9CD203C141402A5AD293C3BABA9",
            INIT_RAM_16 => X"0AD005E832924E92429C091D167806C10041AF32DDE13A669990457D098CC2FE",
            INIT_RAM_17 => X"9A2921ED6AA0CC8387B267B9E7A182720833CEE061E6450C8E4A72E3C087F21A",
            INIT_RAM_18 => X"89A4D43867379AB880C1ACE279E8DA4B3A9063A0B320F65E536B8EAF9CBB9C76",
            INIT_RAM_19 => X"20C76D6362915156A7671331CE657011862E594E46A6D99992E2D640D7668693",
            INIT_RAM_1A => X"3AB1F9007B8A7F2936D16234F9BF9B6BABD48FCE74047C1E738C5B303E815BA7",
            INIT_RAM_1B => X"023170C5DBCC2B6AD72B8E4CCC94DAA079D8BA64E3384337426E7F274CC88A37",
            INIT_RAM_1C => X"144A4566F47B73C95BE6CDB9E664D536762E9224D70F9A5C374B4D1CAB8DF527",
            INIT_RAM_1D => X"7DA5F4A8458A9451315B681ADA9AB0D63218DFB77D3353C32837E954604B9D98",
            INIT_RAM_1E => X"F7D3C6CC8C7841AB49CC538E8A72F2E73C64D2DF3662B19407D7D299CBEDEF3E",
            INIT_RAM_1F => X"77A47C739FF6A22B8B5CDC49E748E9C739BDE6756DB4D22437E74183E12400CB",
            INIT_RAM_20 => X"177AF49DF118FE47ACE3344964FD4ADCFBB543F7729CCB340866D1157B6CCDDB",
            INIT_RAM_21 => X"D6E60DC661155EC9E80F8CEE659F19CC554B2C67C33EDCDA63BAD91B7D1842A7",
            INIT_RAM_22 => X"00FDF3B9B8DE5B76E97F8D32F0F39E4CAC68D9BBB68EA3915F6225F932CAAFDA",
            INIT_RAM_23 => X"441A0CC068A0823F8668A00621B779DE35FEC004050469F34866AEE766743D8C",
            INIT_RAM_24 => X"DA00FADB1D3A630BA18050635DE7DCB13B9B86E0CE6E08DC46331A352F716E3C",
            INIT_RAM_25 => X"A5D31B86A0288D29CE2EAAFF86A6A9F3000082293E6BB54F06698ECCB199973E",
            INIT_RAM_26 => X"D972662C0D31E34E63B31CFC6EB4B35A69B67D85489E62AA99899A94F6800FDB",
            INIT_RAM_27 => X"7FC8531A7A319F3EBFC1383FFCDB0E09BD288288B078B4AD220B6FA934CF6187",
            INIT_RAM_28 => X"96450B74E95A860FF3E434C65F1308F16F92395816B914F0CE870C1323347A4E",
            INIT_RAM_29 => X"7D8C4C59396600DC0C420495A0D987501490002BAD38012E20620D556A230B17",
            INIT_RAM_2A => X"315502751655F60070E6B2C50609369611365AD1E3352327320331A51818030C",
            INIT_RAM_2B => X"AAAC4802B74190FB007C0C0206186AFC1B3A2A46864F26118ED1D03ACB1062B7",
            INIT_RAM_2C => X"E73D9D6D2C265859DB844C2C1952AD10241100174FE0444E6707D80A098D8585",
            INIT_RAM_2D => X"8CF14A288EAE3BFE00FB2DB45080D4A50C58263A3B398DD51AB9CB554ECAA7B2",
            INIT_RAM_2E => X"03AD0025F0D509F63202D877ECD8BF8005451F7BD37367CF0BD9B79850A7D80A",
            INIT_RAM_2F => X"6C60009CA281AEACDC1762945981B869F93D683EAF4AC7EE52412E85B60B91CD",
            INIT_RAM_30 => X"2A191E00538FC8A5004036A959ACB7A463D23E419EA06B744006385455A71250",
            INIT_RAM_31 => X"464C92242004E0AE8518E001D124A7628010115D23C30462FC00A014A1213358",
            INIT_RAM_32 => X"55B555C2278100000A24804D7D98EB98602733818A12094F0B6515022CB40002",
            INIT_RAM_33 => X"4683814663FB910969D1D631A952B381B7F635A33FD38D5CF15DF47D057F7FF5",
            INIT_RAM_34 => X"6A855EC94CFEC4E0172C59A7D054F8F9F4356C312C204E40B05E2059407C8DC8",
            INIT_RAM_35 => X"B38F54EB9091AE3320201EE395AD63902282A031CE3E87CC902954AA515D5D6B",
            INIT_RAM_36 => X"2E5172E82E845070000A846100500E84EA1803B8B07B99E1DC75BE6419674597",
            INIT_RAM_37 => X"A111466C9493A2A7CA2204102414CC798BF0EEC2995A4814580BD07585585ED9",
            INIT_RAM_38 => X"8C2BE27DCB42742742D16797139575DF9649C25019C244097049C2B2DC8D93C4",
            INIT_RAM_39 => X"8C0B50A206C4021E1903C4C176A1A6F73DC560082018912E4371620ACEFC54CB",
            INIT_RAM_3A => X"83B12A14AAB0000B94E92B449483685A51C3067714EA0CC5B1ABA46688C027AB",
            INIT_RAM_3B => X"800000010B5027B80304A59CC71CE149C71CB93D304D209B4C3C61EE98190107",
            INIT_RAM_3C => X"00000000000000000000000000400000856018201DB0516DAAA1FFB5B6DB9241",
            INIT_RAM_3D => X"0A1028440000524A0A4A4A204A5240460800100010540042002064547E060000",
            INIT_RAM_3E => X"8008004042460424402040024A3242124220044022404208520A4A24424A125A",
            INIT_RAM_3F => X"8102080042447C443C0C3C402004FC1838787840407A00707C02487E44487842"
        )
        port map (
            DO => prom_inst_11_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_12: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"A3AE3DB776100108202D7C01D27111171A70BC70EE2CB94289F5EE77F69C7E88",
            INIT_RAM_01 => X"E94F072BF8093090588386DD5449A4199B49C9CA89E96CB003B6D4FEEADB1099",
            INIT_RAM_02 => X"3B401D05F6C97C015DF85D59902EBC0F8FFE050741209036850B689638689B0C",
            INIT_RAM_03 => X"920AC149104E90089A2CF60C1E5D3E2FB862248CD11B593700124C8CAC53E14E",
            INIT_RAM_04 => X"5C6DA844219DC900044879755D55678AC28A24F8D55A006E14698D82D2104BD3",
            INIT_RAM_05 => X"F11BDD946D0844011415415C8AAC0160934C271E30047F2745CD2444BE7A56D7",
            INIT_RAM_06 => X"8528EE337D34514804CEEEE3117C435D6225F37A5774CC56D74DDD3312F5D338",
            INIT_RAM_07 => X"2D24EC5DD2F50F479D513E286F10618467195C6093F2B09BC1D38A88073BB161",
            INIT_RAM_08 => X"566EC5F9B7FFFFF97AAACC90CDE5D7AE3AE14609D432EB4E69F23135FBDE2ADC",
            INIT_RAM_09 => X"CE39FA8ACDC899D73DAECFE29CFFFFFFEAAAAAB93FFF430AFEAAF0FC3F5C5D5D",
            INIT_RAM_0A => X"AD2739A2D1E3D97738FBD598C4048348965FC77A3EDBDDCEB467999D16A961A6",
            INIT_RAM_0B => X"7880187C712481502008C267C6567A3AAE2D910B8CD8A3AC9A7B4EC9C5C01672",
            INIT_RAM_0C => X"7C6DD2FD6605264B58414427C816D9FEEDF8E102BBBDDFB33891C1FBD884A8CA",
            INIT_RAM_0D => X"41E5C4E7022B51115404E2369B959C8C8751C7BFFD7EBCBEFBFDF5E5CF9C0FFB",
            INIT_RAM_0E => X"9095AABEFB5CFB6D196C1B2F0F6202474A0BAA95503531066EEF680444510056",
            INIT_RAM_0F => X"B51F2BD62025C1F26D7FFDBED7B136DB6D56155A49155D3D07FFFED13AD24ED2",
            INIT_RAM_10 => X"998C08889E183BB5C695C59B49623EDDA5B0B4FCDA05D687383A003D8788D138",
            INIT_RAM_11 => X"061D7DB6EFBF493ACBFACCB3EB662B7A12DF7EDB659724986B34444DB706EC5E",
            INIT_RAM_12 => X"F12DCCA5E26219459B7FDF7557DDB2257AB5DE71BFD2DCE22D98F870EB970101",
            INIT_RAM_13 => X"C7A31AC235A1BAF60E5D57FF3FE19767D6DE37FA5BB11273B127706B9AAA5AD2",
            INIT_RAM_14 => X"F3DD75DAD7C5FB55C86205964E5675A3BA639C8E48B30C2200BE1FFBC4816292",
            INIT_RAM_15 => X"D77E723E7FFC9B4E54DD91D1474B93D0D3B6DA30744A9093BA4F74F3DD68EF27",
            INIT_RAM_16 => X"D99FBE660CCE5000F126D175DB427B97B13178CED8EA34BE1FF38D9D37A575B4",
            INIT_RAM_17 => X"866B8AA2AA3C15532240B664C721973C776B772DE8417DE695C5FBDFA1AAAA88",
            INIT_RAM_18 => X"A3BF5CE1A0AA55B5C42B52FF9115EAFA7B2281BA3F60C75786D2AA9621498F34",
            INIT_RAM_19 => X"6D967C9367BCC627DAF781CAB7183F1885A30605C16516CEE725A83E1F1D759E",
            INIT_RAM_1A => X"5E64D734FD979982F28939DEADBE0233E41E478A3BCFB02597249DF5EDA77DFB",
            INIT_RAM_1B => X"05B4029929EA63065338BD4E2F6ABA152B55E20C096FC77B162D3F23CD0129CC",
            INIT_RAM_1C => X"FF898BA36144881500E011C4A304010C05285522D503D6077536AD34786C657C",
            INIT_RAM_1D => X"9C6BC18C0A0D6BAE737FC3EC6294755F0662B154801F3843A3BF79BCDDBA7AB5",
            INIT_RAM_1E => X"15AA76E6BE3E3DD42D65C52F7CBABDFDCD7C71F4CF11D5764F14CCCAB5ABAAD9",
            INIT_RAM_1F => X"9FA000000A6E7EC3C4A02E3447D90955FE5A01108A514257F8D11D5549856D95",
            INIT_RAM_20 => X"A3AE3DB776100108202D7C01D27111171A70BC70EE2CB94289F5EE77F69C7E88",
            INIT_RAM_21 => X"E94F072BF8093090588386DD5449A4199B49C9CA89E96CB003B6D4FEEADB1099",
            INIT_RAM_22 => X"3B401D05F6C97C015DF85D59902EBC0F8FFE050741209036850B689638689B0C",
            INIT_RAM_23 => X"920AC149104E90089A2CF60C1E5D3E2FB862248CD11B593700124C8CAC53E14E",
            INIT_RAM_24 => X"5C6DA844219DC900044879755D55678AC28A24F8D55A006E14698D82D2104BD3",
            INIT_RAM_25 => X"F11BDD946D0844011415415C8AAC0160934C271E30047F2745CD2444BE7A56D7",
            INIT_RAM_26 => X"8528EE337D34514804CEEEE3117C435D6225F37A5774CC56D74DDD3312F5D338",
            INIT_RAM_27 => X"2D24EC5DD2F50F479D513E286F10618467195C6093F2B09BC1D38A88073BB161",
            INIT_RAM_28 => X"566EC5F9B7FFFFF97AAACC90CDE5D7AE3AE14609D432EB4E69F23135FBDE2ADC",
            INIT_RAM_29 => X"CE39FA8ACDC899D73DAECFE29CFFFFFFEAAAAAB93FFF430AFEAAF0FC3F5C5D5D",
            INIT_RAM_2A => X"AD2739A2D1E3D97738FBD598C4048348965FC77A3EDBDDCEB467999D16A961A6",
            INIT_RAM_2B => X"7880187C712481502008C267C6567A3AAE2D910B8CD8A3AC9A7B4EC9C5C01672",
            INIT_RAM_2C => X"7C6DD2FD6605264B58414427C816D9FEEDF8E102BBBDDFB33891C1FBD884A8CA",
            INIT_RAM_2D => X"41E5C4E7022B51115404E2369B959C8C8751C7BFFD7EBCBEFBFDF5E5CF9C0FFB",
            INIT_RAM_2E => X"9095AABEFB5CFB6D196C1B2F0F6202474A0BAA95503531066EEF680444510056",
            INIT_RAM_2F => X"B51F2BD62025C1F26D7FFDBED7B136DB6D56155A49155D3D07FFFED13AD24ED2",
            INIT_RAM_30 => X"998C08889E183BB5C695C59B49623EDDA5B0B4FCDA05D687383A003D8788D138",
            INIT_RAM_31 => X"061D7DB6EFBF493ACBFACCB3EB662B7A12DF7EDB659724986B34444DB706EC5E",
            INIT_RAM_32 => X"F12DCCA5E26219459B7FDF7557DDB2257AB5DE71BFD2DCE22D98F870EB970101",
            INIT_RAM_33 => X"C7A31AC235A1BAF60E5D57FF3FE19767D6DE37FA5BB11273B127706B9AAA5AD2",
            INIT_RAM_34 => X"F3DD75DAD7C5FB55C86205964E5675A3BA639C8E48B30C2200BE1FFBC4816292",
            INIT_RAM_35 => X"D77E723E7FFC9B4E54DD91D1474B93D0D3B6DA30744A9093BA4F74F3DD68EF27",
            INIT_RAM_36 => X"D99FBE660CCE5000F126D175DB427B97B13178CED8EA34BE1FF38D9D37A575B4",
            INIT_RAM_37 => X"866B8AA2AA3C15532240B664C721973C776B772DE8417DE695C5FBDFA1AAAA88",
            INIT_RAM_38 => X"A3BF5CE1A0AA55B5C42B52FF9115EAFA7B2281BA3F60C75786D2AA9621498F34",
            INIT_RAM_39 => X"6D967C9367BCC627DAF781CAB7183F1885A30605C16516CEE725A83E1F1D759E",
            INIT_RAM_3A => X"5E64D734FD979982F28939DEADBE0233E41E478A3BCFB02597249DF5EDA77DFB",
            INIT_RAM_3B => X"05B4029929EA63065338BD4E2F6ABA152B55E20C096FC77B162D3F23CD0129CC",
            INIT_RAM_3C => X"FF898BA36144881500E011C4A304010C05285522D503D6077536AD34786C657C",
            INIT_RAM_3D => X"9C6BC18C0A0D6BAE737FC3EC6294755F0662B154801F3843A3BF79BCDDBA7AB5",
            INIT_RAM_3E => X"15AA76E6BE3E3DD42D65C52F7CBABDFDCD7C71F4CF11D5764F14CCCAB5ABAAD9",
            INIT_RAM_3F => X"9FA000000A6E7EC3C4A02E3447D90955FE5A01108A514257F8D11D5549856D95"
        )
        port map (
            DO => prom_inst_12_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_13: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"A3AE3DB776100108202D7C01D27111171A70BC70EE2CB94289F5EE77F69C7E88",
            INIT_RAM_01 => X"E94F072BF8093090588386DD5449A4199B49C9CA89E96CB003B6D4FEEADB1099",
            INIT_RAM_02 => X"3B401D05F6C97C015DF85D59902EBC0F8FFE050741209036850B689638689B0C",
            INIT_RAM_03 => X"920AC149104E90089A2CF60C1E5D3E2FB862248CD11B593700124C8CAC53E14E",
            INIT_RAM_04 => X"5C6DA844219DC900044879755D55678AC28A24F8D55A006E14698D82D2104BD3",
            INIT_RAM_05 => X"F11BDD946D0844011415415C8AAC0160934C271E30047F2745CD2444BE7A56D7",
            INIT_RAM_06 => X"8528EE337D34514804CEEEE3117C435D6225F37A5774CC56D74DDD3312F5D338",
            INIT_RAM_07 => X"2D24EC5DD2F50F479D513E286F10618467195C6093F2B09BC1D38A88073BB161",
            INIT_RAM_08 => X"566EC5F9B7FFFFF97AAACC90CDE5D7AE3AE14609D432EB4E69F23135FBDE2ADC",
            INIT_RAM_09 => X"CE39FA8ACDC899D73DAECFE29CFFFFFFEAAAAAB93FFF430AFEAAF0FC3F5C5D5D",
            INIT_RAM_0A => X"AD2739A2D1E3D97738FBD598C4048348965FC77A3EDBDDCEB467999D16A961A6",
            INIT_RAM_0B => X"7880187C712481502008C267C6567A3AAE2D910B8CD8A3AC9A7B4EC9C5C01672",
            INIT_RAM_0C => X"7C6DD2FD6605264B58414427C816D9FEEDF8E102BBBDDFB33891C1FBD884A8CA",
            INIT_RAM_0D => X"41E5C4E7022B51115404E2369B959C8C8751C7BFFD7EBCBEFBFDF5E5CF9C0FFB",
            INIT_RAM_0E => X"9095AABEFB5CFB6D196C1B2F0F6202474A0BAA95503531066EEF680444510056",
            INIT_RAM_0F => X"B51F2BD62025C1F26D7FFDBED7B136DB6D56155A49155D3D07FFFED13AD24ED2",
            INIT_RAM_10 => X"998C08889E183BB5C695C59B49623EDDA5B0B4FCDA05D687383A003D8788D138",
            INIT_RAM_11 => X"061D7DB6EFBF493ACBFACCB3EB662B7A12DF7EDB659724986B34444DB706EC5E",
            INIT_RAM_12 => X"F12DCCA5E26219459B7FDF7557DDB2257AB5DE71BFD2DCE22D98F870EB970101",
            INIT_RAM_13 => X"C7A31AC235A1BAF60E5D57FF3FE19767D6DE37FA5BB11273B127706B9AAA5AD2",
            INIT_RAM_14 => X"F3DD75DAD7C5FB55C86205964E5675A3BA639C8E48B30C2200BE1FFBC4816292",
            INIT_RAM_15 => X"D77E723E7FFC9B4E54DD91D1474B93D0D3B6DA30744A9093BA4F74F3DD68EF27",
            INIT_RAM_16 => X"D99FBE660CCE5000F126D175DB427B97B13178CED8EA34BE1FF38D9D37A575B4",
            INIT_RAM_17 => X"866B8AA2AA3C15532240B664C721973C776B772DE8417DE695C5FBDFA1AAAA88",
            INIT_RAM_18 => X"A3BF5CE1A0AA55B5C42B52FF9115EAFA7B2281BA3F60C75786D2AA9621498F34",
            INIT_RAM_19 => X"6D967C9367BCC627DAF781CAB7183F1885A30605C16516CEE725A83E1F1D759E",
            INIT_RAM_1A => X"5E64D734FD979982F28939DEADBE0233E41E478A3BCFB02597249DF5EDA77DFB",
            INIT_RAM_1B => X"05B4029929EA63065338BD4E2F6ABA152B55E20C096FC77B162D3F23CD0129CC",
            INIT_RAM_1C => X"FF898BA36144881500E011C4A304010C05285522D503D6077536AD34786C657C",
            INIT_RAM_1D => X"9C6BC18C0A0D6BAE737FC3EC6294755F0662B154801F3843A3BF79BCDDBA7AB5",
            INIT_RAM_1E => X"15AA76E6BE3E3DD42D65C52F7CBABDFDCD7C71F4CF11D5764F14CCCAB5ABAAD9",
            INIT_RAM_1F => X"9FA000000A6E7EC3C4A02E3447D90955FE5A01108A514257F8D11D5549856D95",
            INIT_RAM_20 => X"A3AE3DB776100108202D7C01D27111171A70BC70EE2CB94289F5EE77F69C7E88",
            INIT_RAM_21 => X"E94F072BF8093090588386DD5449A4199B49C9CA89E96CB003B6D4FEEADB1099",
            INIT_RAM_22 => X"3B401D05F6C97C015DF85D59902EBC0F8FFE050741209036850B689638689B0C",
            INIT_RAM_23 => X"920AC149104E90089A2CF60C1E5D3E2FB862248CD11B593700124C8CAC53E14E",
            INIT_RAM_24 => X"5C6DA844219DC900044879755D55678AC28A24F8D55A006E14698D82D2104BD3",
            INIT_RAM_25 => X"F11BDD946D0844011415415C8AAC0160934C271E30047F2745CD2444BE7A56D7",
            INIT_RAM_26 => X"8528EE337D34514804CEEEE3117C435D6225F37A5774CC56D74DDD3312F5D338",
            INIT_RAM_27 => X"2D24EC5DD2F50F479D513E286F10618467195C6093F2B09BC1D38A88073BB161",
            INIT_RAM_28 => X"566EC5F9B7FFFFF97AAACC90CDE5D7AE3AE14609D432EB4E69F23135FBDE2ADC",
            INIT_RAM_29 => X"CE39FA8ACDC899D73DAECFE29CFFFFFFEAAAAAB93FFF430AFEAAF0FC3F5C5D5D",
            INIT_RAM_2A => X"AD2739A2D1E3D97738FBD598C4048348965FC77A3EDBDDCEB467999D16A961A6",
            INIT_RAM_2B => X"7880187C712481502008C267C6567A3AAE2D910B8CD8A3AC9A7B4EC9C5C01672",
            INIT_RAM_2C => X"7C6DD2FD6605264B58414427C816D9FEEDF8E102BBBDDFB33891C1FBD884A8CA",
            INIT_RAM_2D => X"41E5C4E7022B51115404E2369B959C8C8751C7BFFD7EBCBEFBFDF5E5CF9C0FFB",
            INIT_RAM_2E => X"9095AABEFB5CFB6D196C1B2F0F6202474A0BAA95503531066EEF680444510056",
            INIT_RAM_2F => X"B51F2BD62025C1F26D7FFDBED7B136DB6D56155A49155D3D07FFFED13AD24ED2",
            INIT_RAM_30 => X"998C08889E183BB5C695C59B49623EDDA5B0B4FCDA05D687383A003D8788D138",
            INIT_RAM_31 => X"061D7DB6EFBF493ACBFACCB3EB662B7A12DF7EDB659724986B34444DB706EC5E",
            INIT_RAM_32 => X"F12DCCA5E26219459B7FDF7557DDB2257AB5DE71BFD2DCE22D98F870EB970101",
            INIT_RAM_33 => X"C7A31AC235A1BAF60E5D57FF3FE19767D6DE37FA5BB11273B127706B9AAA5AD2",
            INIT_RAM_34 => X"F3DD75DAD7C5FB55C86205964E5675A3BA639C8E48B30C2200BE1FFBC4816292",
            INIT_RAM_35 => X"D77E723E7FFC9B4E54DD91D1474B93D0D3B6DA30744A9093BA4F74F3DD68EF27",
            INIT_RAM_36 => X"D99FBE660CCE5000F126D175DB427B97B13178CED8EA34BE1FF38D9D37A575B4",
            INIT_RAM_37 => X"866B8AA2AA3C15532240B664C721973C776B772DE8417DE695C5FBDFA1AAAA88",
            INIT_RAM_38 => X"A3BF5CE1A0AA55B5C42B52FF9115EAFA7B2281BA3F60C75786D2AA9621498F34",
            INIT_RAM_39 => X"6D967C9367BCC627DAF781CAB7183F1885A30605C16516CEE725A83E1F1D759E",
            INIT_RAM_3A => X"5E64D734FD979982F28939DEADBE0233E41E478A3BCFB02597249DF5EDA77DFB",
            INIT_RAM_3B => X"05B4029929EA63065338BD4E2F6ABA152B55E20C096FC77B162D3F23CD0129CC",
            INIT_RAM_3C => X"FF898BA36144881500E011C4A304010C05285522D503D6077536AD34786C657C",
            INIT_RAM_3D => X"9C6BC18C0A0D6BAE737FC3EC6294755F0662B154801F3843A3BF79BCDDBA7AB5",
            INIT_RAM_3E => X"15AA76E6BE3E3DD42D65C52F7CBABDFDCD7C71F4CF11D5764F14CCCAB5ABAAD9",
            INIT_RAM_3F => X"9FA000000A6E7EC3C4A02E3447D90955FE5A01108A514257F8D11D5549856D95"
        )
        port map (
            DO => prom_inst_13_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_14: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"7EF77AB52F01EF7FF323C9F5287DAEBACF8FC472607DBA848425C4090B09013C",
            INIT_RAM_01 => X"02C344D85A48A3249394F5AC934726B4D591CAAB3B5DB529ED77B22422D829B2",
            INIT_RAM_02 => X"7F5AC3A9F0DF87EF2E6537D65EF7B6F2D61962A74ECD62C5E336A8A9C2676DC9",
            INIT_RAM_03 => X"6EA0A65EF790517FCF3BF7C7859D49E588FE5FB306243EDC5D596997B0D645BD",
            INIT_RAM_04 => X"41998C465331908C20D64088C620110000001953FE882B83ACFA8DF9E2A5F777",
            INIT_RAM_05 => X"4A1EB6CFFFE773E7DFF9C0040E10AD08A5005632313588448446982A8CCC0066",
            INIT_RAM_06 => X"779FFE342C44241118E9E4538A31BB3773DBA67F1A6BADF6F261DB2BFE37834F",
            INIT_RAM_07 => X"E8BACAFAE413AB0456AF49CE172F1071E1E7F4D0B8C168F59CC37630F4B99A3F",
            INIT_RAM_08 => X"2FD4E81379CDAC4A870CFBB26BB54875D77B1D8EEAEB9A66FDB99DE6E236D42E",
            INIT_RAM_09 => X"83032916F692AA32AA23333E9485A80A3554705242808F0A9C7A5617969F13CF",
            INIT_RAM_0A => X"8F8B149733D523AF47F6DF4DAAFD3F5BF242E8C4B26423FFF243F7EF8A9A3B28",
            INIT_RAM_0B => X"D3DBE37192D5DA0E63AAF7F24B3F6DBF6792DA7BFEF081395C287B0591E88D25",
            INIT_RAM_0C => X"7E67E637FF7DF7C4FE737F3663FE71FD2AA1346D1574C071BE3F64DD54C75731",
            INIT_RAM_0D => X"0762FCBFFAAAAF0AC82C192D0C14EF1F3FBC3350E85A8FF6EDA50516BCEBF9DF",
            INIT_RAM_0E => X"DE3EF2C425F72CEFD375BFDDDBE5F979CFFA7EF4CDB8202CF9F71E27FA92CA70",
            INIT_RAM_0F => X"BC2A2E535906BBF727E98A064DFD1CC215BF37D94BAB6B7EF6F6F4F4F6F72507",
            INIT_RAM_10 => X"415541114044101500116BEBFBFF37D94BA7FA374ED77617A8359050BF20BE94",
            INIT_RAM_11 => X"79B1E6BE008ABEFAE857F7ECA59272AACB24D555550001554055054145104451",
            INIT_RAM_12 => X"5A35FC0BDF99097745A3EC76FDAD7CDB54D7E8D37150675D0FD7CBE3969C4F8C",
            INIT_RAM_13 => X"5B628E5986455437CE610D055A955BFF54DDE2CF07DB1B77EF96002E17FC7775",
            INIT_RAM_14 => X"E36FB4955BE8D6FB7DA6B5FDEB599B6FB46AD36DAD5A6AD5ADED1FBA60A6D1B1",
            INIT_RAM_15 => X"18ECEDF2F4A54925E22B69B208060F42C1F59A2B3B6131F783F64E8ABB35F6AB",
            INIT_RAM_16 => X"8A977F82E8DD9721358D8910C5EC3D88CE864430A41F60633194C23BEC7029D0",
            INIT_RAM_17 => X"AF59A954553EE6D6767D9F7DE406E1A03AFD25E7F8BBED36BA5BCAAFAAD0A76B",
            INIT_RAM_18 => X"5F889B26EBE9BAF13310EF167F1AD5B194C58DDAD90EF6FF667BBCD34EB92651",
            INIT_RAM_19 => X"D5375EBF87CDE595FDDEFB60000B7BD62B9D5B07370B2AFB59BD6574EFEF7DFB",
            INIT_RAM_1A => X"736DB066EB1A38228B3BAC6239EDB33636FC68AD2C55A2C498ACA2FBFEB1ED17",
            INIT_RAM_1B => X"E92D317BADF77C55A5DD3B7B7E6DDE5948AA6768EA3CC84C9003EB391CD68FC4",
            INIT_RAM_1C => X"7DDE71ADB679E79AA165F0F936E2C6013ECBB90DD6DB4EEB54BA775FA698BDD4",
            INIT_RAM_1D => X"975C380628580C094BD85DB7CCBB6FFAD5BD96C39D753CF3CCAFB1695ED4DF27",
            INIT_RAM_1E => X"76CF15E24E87743358AB8A9358AB5975C018A1700600484AC2B4335CA9358EB5",
            INIT_RAM_1F => X"4611E7BEEDFCEFBC5BFC49C7FAD5BDF7FADBEF32FEBE6E36F37E6E73EC49D0E8",
            INIT_RAM_20 => X"28E49593A85722FB048B0AC493449976DA25EF78AA5F7D0D78FB4AD8FB61E91C",
            INIT_RAM_21 => X"E6F9DEDAC4B36A6BEED5D24D23CB9DFCA55AB9BCE02699B5541FF8019A48F8A7",
            INIT_RAM_22 => X"FD87F9A8BBBCE8DFFDD4A47DE5DBE5F315EA4675C54EAC43ED285C9BC1D9F36E",
            INIT_RAM_23 => X"CCB01672062A1D8EEE03804F8705B33AB8F201AC7D9183C959A5B7A33A5CD736",
            INIT_RAM_24 => X"1B761EFA5BD298A5BAA8A71EEEF443B951585DDF7E30B222222236297A88C2F6",
            INIT_RAM_25 => X"F8EF1F7E65B36862F88205B35BC338720B0750C3FD74B6FB6D192947D0C75347",
            INIT_RAM_26 => X"06991FC69FFBBFFBACD687E37C995D9503803DB3E6F5AE0BDB4FBF017D1EBC9E",
            INIT_RAM_27 => X"5220019249CB019900A21272D2400004249108182089268805B8A718FF4D9F74",
            INIT_RAM_28 => X"7C4D94CB0000B86FC2AC13E1E19FD7D80BEEE9D5D80F18CAB4EAAF0EEF764400",
            INIT_RAM_29 => X"E5155F7FB3F877DA7EAF7C3BED3E8F7C4307FCEFFB8D417D5BFF76AFF4F9BD4E",
            INIT_RAM_2A => X"D59EEFFCFFE79DF515F9CAFA8EFD97ECFF295F0AB1D7EF39C3AC55F70A054502",
            INIT_RAM_2B => X"F75E72524A49E8A8A6EE0A8C79E09E1DBC9FCBBFA5E8CF03C542B66F0942BD3A",
            INIT_RAM_2C => X"88F255A7BF5ED75AE0208122CCC1660DF6E0DF9E5A704E8BC608B6DF5B8FB9F1",
            INIT_RAM_2D => X"B8AA7291C7DE2A9CB86B447E6A9CED9055AF92322BCAB7C31E42F318F69456DA",
            INIT_RAM_2E => X"0000420E8B86665712B8BA6EC34CC42DE45A31E5E0C3B479A661DA6704CBFE49",
            INIT_RAM_2F => X"6172A5E3E4A53CE914C8E0347F9F093892222569201540A18708F6E2BC088000",
            INIT_RAM_30 => X"CA81AD206010B0AFA14E55DBD830CEE549E71D2BB6D6F3045507C944B8DDE1C5",
            INIT_RAM_31 => X"ECC9502A82A97014C712207F38AF70B53C48374851A0BCA0906680382215449C",
            INIT_RAM_32 => X"DBC0F04080924924E346B1FBC863D96CD8238240323F902C3ED2C6CB2280E034",
            INIT_RAM_33 => X"04CFC93502265E62C700A3420D08119114CAB0982626262313456C8B92DDFD6A",
            INIT_RAM_34 => X"E82D026BE3443471B8E8966497FB70123CE30E38CCA5837B06E3DC5E3B6166D8",
            INIT_RAM_35 => X"187C36676672993B2032602AA80D682D90E9028E6E540BD2F540FD8976C26E64",
            INIT_RAM_36 => X"31562C8A0298E0551144E6BA2A32CFFE5A472ECC616843D08B0C08F0C08E0C09",
            INIT_RAM_37 => X"020008859ED08271F5A7C5F5B3C86B61B434718E8D45D5BA16ED4EC1C177870F",
            INIT_RAM_38 => X"66220EDD1456AFEF7BD21EC436ED6DC11ECC1509282B1A883265468200001FE2",
            INIT_RAM_39 => X"DF0E9550E2A7FF7512378BA7962B21F4DBBE287FA9376D4E7888EE7DAB070CD3",
            INIT_RAM_3A => X"C00826E25FBBF1944E8E127471A5B476A05030BF80C06B75CED132ABC2EAECF6",
            INIT_RAM_3B => X"2A126B12593BBAFFF8B4FFFA8B9BD23BC1223EFBFAB7C06512DCAB9FC492107B",
            INIT_RAM_3C => X"D91D7FC55C62ECFE2748DF8B84F1A6E917B20CADE97751CCECDAAA4F7B8BDBE8",
            INIT_RAM_3D => X"9CB9EE85D6669AEDB2AED69EB348ADC14EC1C66C03BFE9F665298CFE1DF7C8FD",
            INIT_RAM_3E => X"2FE17F2AEBF2C472EFE10846BD7DEFBE359E237577995DA6E6B3DB5FC3B5825B",
            INIT_RAM_3F => X"30016EF3219421AE121CFCDCF4D4DC4BC66B1F7347A4A020BEB2BEC56CEFDBD6"
        )
        port map (
            DO => prom_inst_14_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_2,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_15: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"CC8070206B8245AC240020752EBC2BEF3E748D3F8F361C239C4AFAE93FF8775A",
            INIT_RAM_01 => X"00812F408CC6501331852531B04480021D9220D4903A41404312032840153FE9",
            INIT_RAM_02 => X"B383E6E7C3B310E1F7FF595C5DF6F0E9A9FFFBE16D3FFBE82C1E0051F1E060D5",
            INIT_RAM_03 => X"C1FFFB3487617BE24FD79501DE05F1A341B89EC82FD5702597FD866639C0DE08",
            INIT_RAM_04 => X"47A8EA413A2DCF0BFA8EEC2318DBF3C4711871B3BC0404EC45252A485234A663",
            INIT_RAM_05 => X"1D2FCA8DCB43C5356BAE638588C302868CE1161CACADFEF7696F8C3AA82EC16F",
            INIT_RAM_06 => X"FF4DEBFBDEB376DF68D5EEDB5EB4D5AB5B39745D76CD8ADC59CB30C8AA33E155",
            INIT_RAM_07 => X"06ABC52D5DBEF57EEB3311A9D85D253B44E250E1566BED57C6DFEB2ABFD1ADF6",
            INIT_RAM_08 => X"D7D77EF5E2C6D7220BE64B3C6E9EF22AFDFCC8005C2FFFFA3AB9AD1ADFC0AFE7",
            INIT_RAM_09 => X"DCD4560015805B13AC0290001EF826137E4EB867C828D9777FFF47B6903008DD",
            INIT_RAM_0A => X"1C9DCD8EBB9D36AF570CF25CDD16F645D1DE9F9EE575E2A2B91D5659FC131CE3",
            INIT_RAM_0B => X"CF133BF47B9D3DA46DD6DBF3A8ADCDD3DF1176D2FE1B447DFC65E1DD7BF3BE5E",
            INIT_RAM_0C => X"F0A09C47F23F20FE2ACFF5FD3ABE6167E5FD36E1D9735BBD5375C1F79BD0424E",
            INIT_RAM_0D => X"3497229CB9044B6E7A7861A04A712AAF29EFBD393727F1F3FC2AB1E6CF571457",
            INIT_RAM_0E => X"A8BCDC266655185CC45008B39EFD1FA6E9F5E816114F93E1E7A2A27C72C7349F",
            INIT_RAM_0F => X"FD5CB07B6C729B510A78BEC5F7C7A1E7809F1976D0DD3615C1D27D2DF596BFE7",
            INIT_RAM_10 => X"63B065F7D671322D6BFB2B8759433929CEC27E3FD7741292A4A5AF02703CF4E3",
            INIT_RAM_11 => X"DDB3A42AC80797FDEF4DE3EEF7ED8C7307E4CE6A6317F7BF25D077BBF03AEA33",
            INIT_RAM_12 => X"59BD7F8DE9FBF27A65DE5245BEBC7DAA0A70DB7240B0D136169D77D649A39EB4",
            INIT_RAM_13 => X"21A40982C046D22C10146484345CAF7BC828BFE79DFBEFC4B1CBF660C487EBB7",
            INIT_RAM_14 => X"CCCA0665222D038CC873351A21B23939A98CC08803282189C8440D40CD404624",
            INIT_RAM_15 => X"9CD4E55E6CB00410842B02A7FD105706DF9E2A1FA025005632A0CC080400D280",
            INIT_RAM_16 => X"130E0174D4FB44B2C0D7A907702A748D0BA50F8FA5437ACD3B343C35039F44D1",
            INIT_RAM_17 => X"8AB3B7FDEE7B9CC735FCCE93E3AC1AAAA691AD6350E57F1F5773302B6072C63D",
            INIT_RAM_18 => X"F7F22D2FE1509BDF80E6DD7B7175B71C6531C3A86BE9F1D7A6AFD5FFB7A37A60",
            INIT_RAM_19 => X"7CA976FE488D1069D687A6F1D68A70F37CAAA367A74CBB73D3A6FFB4B1E8D4B7",
            INIT_RAM_1A => X"681A00AF8D864D8BB6D2A0916C8A9B250A76B8A977F82E8FDFBE68F8E0F8DF23",
            INIT_RAM_1B => X"BFF05FBD6AD8CA62C6CBE43BDBFD99E8EB6DD724D235FBEA9FE7D6767D811C40",
            INIT_RAM_1C => X"AF72F66DC666B39A6D66FD958ED9BC6D758D5EC24DFEBA64871D6B86D37DF1DF",
            INIT_RAM_1D => X"FBB9EB400590D7F939FF5A70A29817DC2CC29B679B2D7146BD21D47EF06F7D5E",
            INIT_RAM_1E => X"B4B15EB89456517DFF58F68BDADB95B5F764CBE7E7C7E7DF0CADB8FFD8F9A72B",
            INIT_RAM_1F => X"7BBD7F79FFE0AB8FC33758D1C1145DDD6311CF69FFFDF62EDD236FC6A0358FA2",
            INIT_RAM_20 => X"26FAFE3BE30DFAF7B9E7A5FFE4797314DAA1C1529CDBFFE9D94EB11A9F68D4DF",
            INIT_RAM_21 => X"A1FF3BE5E159FFDDEB2FBECAEB87BBCC5FCF6E23D77E4DD4C9DEBC93C10F6363",
            INIT_RAM_22 => X"2175C7B89C48CCC916D46F9315DFDECBE43E5F03D7D27F97E09E4700AA694552",
            INIT_RAM_23 => X"768008002000002624793100811F43BC315A6004052671392B47FEB7F5DC90E6",
            INIT_RAM_24 => X"8ED67F67AA66B0674CD240410F613700B8DFE7F8837F88FF4520002E4BFD7FA2",
            INIT_RAM_25 => X"7941B61372AC884EE60A372057B59CF990A6020B875C06E7C53BDF9A91F8F058",
            INIT_RAM_26 => X"8CA3CE9F24BEFA9E2BB9D89B423C327C8E050114401A63BDCD2054E166C0005F",
            INIT_RAM_27 => X"420539B476E305B8200E47DFAAE8D5D1D0724DCC3FD72C4F8DE54622A1DD1BA7",
            INIT_RAM_28 => X"EF3142B9927BEAF99BCFB066319F5BDF2EFFB11686607A73BE9CB85CF6EC52D0",
            INIT_RAM_29 => X"E3BE607B3FAC5DD39FB436C5BB7926D7FFF03EF787FF563C3FEF787919A8383D",
            INIT_RAM_2A => X"EB9963425C951C00298F26A884C3AEF0DBF539D04E867EB6FB957E817C230DFE",
            INIT_RAM_2B => X"3DDBF48E39F1AE9FC0A7CAC2B4515882877D84D415C7A00D91E87F57E95B60EF",
            INIT_RAM_2C => X"86E8AEC1EE37F6F5FFD77F204F5EBFDA614C41C1F85C32FFB05F2881BF7EB1D7",
            INIT_RAM_2D => X"60BE688D11B16D7936F4B55E0E301BAD6A96802B5719271D55D5E93FEE5335EF",
            INIT_RAM_2E => X"04FF86DDFE9FCBD3DC2A4967F492CDD5A8FFBD98573036C583F9D6D6A6138C03",
            INIT_RAM_2F => X"CE21FFE0D222852612C7A87E8DFE961BD8CF052D4757559DF3ED2417472384AF",
            INIT_RAM_30 => X"35995E3ADF9E07EB861E3035B1EF3EF935DAFFFA1F94FDCA5B833F14101BE318",
            INIT_RAM_31 => X"896B7EB5FD69B679669CBA00AA9A431956A3CE676A9D7B50D84F3FFFFFC4AAF7",
            INIT_RAM_32 => X"AA8AAA32A2C38012BFEB492278CD27651FD91BDE452EEF053E0D2912A0D49D9A",
            INIT_RAM_33 => X"C165510222E12BABC9B940EB70182EDBEEF007365AA980A2002829A05282A2AA",
            INIT_RAM_34 => X"F70811E17D8C73F1D9BEF7F7E82EFAE6C2D2DB2126004D81CA67DACC344F6458",
            INIT_RAM_35 => X"776B42A5FE80BB5AAA2A550A58904A1C6DC992952AB4532C6CB2F975BC101356",
            INIT_RAM_36 => X"4B7AE34419240F3C0170E001D6CE75F0475D5A8A9012B9BD97153AB038EF6187",
            INIT_RAM_37 => X"812017671773A9EE08641F818054455F0BABE232D2AA00081423C0BCCE1E642C",
            INIT_RAM_38 => X"B4A728E3A780E88E8A333EFF77B3F75DD75370020203478F160F42F9A061FE44",
            INIT_RAM_39 => X"B1D336B62293FF5CBBEE347FBBF8EF6BF394BB6DBDDECE9C3FDDE42969D88FED",
            INIT_RAM_3A => X"9559B18B257000031ED659F13ED53E8F9B9F2F6623EE2875FBD95BED308D5057",
            INIT_RAM_3B => X"800000012A022D0E60C9CC6E8469ED13069CBC7878F870A2183FBE417F1DC1DB",
            INIT_RAM_3C => X"000000000000000000000000002473989D7348225CA8053DA57353A59FFF9249",
            INIT_RAM_3D => X"522828280000524A124A4A7E4A527E4A106010607C38003C025408FE24000000",
            INIT_RAM_3E => X"800400207E4A0818204040024A1262124210084014407E08520A4A42424A1256",
            INIT_RAM_3F => X"A504087E764CA02840304044540424244404044024804008A40A54484448544A"
        )
        port map (
            DO => prom_inst_15_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_16: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"97E42BA702155AF7AB422B5B647561935CD2B6357F49C99DC983C8F6D01A728B",
            INIT_RAM_01 => X"1250010D180454827A0E040040692415D222BA8E29DCEF710B77D8FC4B52B025",
            INIT_RAM_02 => X"B653590C7D810C15C2857B460280048007FE0801004D2BA423904104201D5215",
            INIT_RAM_03 => X"0568C11050163AAA612C780C2E983DC490024315217110A456BC353502D20A08",
            INIT_RAM_04 => X"28560460E9245100030C0DC251A4C1D402CC614261A2115B000411D1DA015DD0",
            INIT_RAM_05 => X"E150BB2941090150451488BC8FC501063AEC015CFC76D56C55E4A71632326293",
            INIT_RAM_06 => X"01040000259B5A62A9ACCCDE0502A0A018B190726B649948C64AD92658C1922A",
            INIT_RAM_07 => X"C848D5818383860F806126680D9037AC441004840AD4310760819046A55808E5",
            INIT_RAM_08 => X"20D183053A15555331409B059BFB6410410CC8ABD6B494944DE0A7830B150AAF",
            INIT_RAM_09 => X"123A1485B9890197750FD6AA9E0400000010000415551504545041A86AC2EB20",
            INIT_RAM_0A => X"205B3D9D0297823E748119980000820916545050BF77E6605547AECF964EE102",
            INIT_RAM_0B => X"3D007F8C502301204003B2E4508E702C2EA81209D6FABAAFA23FC2D9C95F2AE5",
            INIT_RAM_0C => X"3C6FF4EDD615D01204B26DEFD363924001E870257A3C895F91F1A3E1E55A3320",
            INIT_RAM_0D => X"AE5555B502A7F5854894C0A11594BD3E8D70C58B767050998C8DBCE48B9D1FCB",
            INIT_RAM_0E => X"E0DFC3D5EFE9CFFF43B09D340628202CE2031554847244445554D6ABEAABEBEE",
            INIT_RAM_0F => X"3D0C20468221A9E6FFEA9996ADAEC136D8824A8EDB4001A80EAAA8636C76D860",
            INIT_RAM_10 => X"CEAF2A21C40C3BCE12C191C6FFDE3D7A86600ACE99D18905A18C846FA18BAF48",
            INIT_RAM_11 => X"1CE8F7FFADFDFFEB7F376897C02D0168425BFBFFD6FEFFF48FE5908A6E533935",
            INIT_RAM_12 => X"F0A07071F12B76DF4318E73EA199B60E7ECC21D69B8AE180C8AAD020EC484611",
            INIT_RAM_13 => X"037E88EE753608120730E5543EA759DD9DB2D3715C52E9CC86A63200E5503CFA",
            INIT_RAM_14 => X"6DA7FDA97D80A29960EC0F8BE70DDA56ECA30C00706904C1348C27B28A214C02",
            INIT_RAM_15 => X"5F1F37CC47502BFDC6015E1EDDA326A6C51CF3C1F90BF3319964D3F7F3F9280F",
            INIT_RAM_16 => X"9AB36CE939D8C505D7926380E1284510EF807B2E70E3CE2DBA8577FBC238DDAB",
            INIT_RAM_17 => X"4E8A1C5554D14A124FD73F32692136B898DB3C3356D3748EE1F3EC99712C32AF",
            INIT_RAM_18 => X"C6CC08D082742C7B9C8A4186E00BAEDDA466C3924D365936D966003EC0D70698",
            INIT_RAM_19 => X"DB5BDBFED6111060952622150248737130E9AD230A82E32DAC06101D3B4B428E",
            INIT_RAM_1A => X"9EEA7DEDDD27BA52A5212180A0814001841C475661CE2084B66DB12D9B6C4B66",
            INIT_RAM_1B => X"4574449909AA2281574ABDC2AF4018098038110245A0D7EC78097700D04E83A4",
            INIT_RAM_1C => X"CCA8CEF241448805A0E251C4A504250C150615269527B51B63348F117E2C6C7C",
            INIT_RAM_1D => X"9837615FEC2937278B31E19B3B14642A1D68E50D881930D387DF99CCCC9F9E61",
            INIT_RAM_1E => X"139ACE6EBC36ACB8AD93EA23D4387D9CDD786BDA6D4ED82E049AAAAD89DCCDE5",
            INIT_RAM_1F => X"72A0000002E29E9405902E12574985A854381210B4A152970A521A861B83A528",
            INIT_RAM_20 => X"97E42BA702155AF7AB422B5B647561935CD2B6357F49C99DC983C8F6D01A728B",
            INIT_RAM_21 => X"1250010D180454827A0E040040692415D222BA8E29DCEF710B77D8FC4B52B025",
            INIT_RAM_22 => X"B653590C7D810C15C2857B460280048007FE0801004D2BA423904104201D5215",
            INIT_RAM_23 => X"0568C11050163AAA612C780C2E983DC490024315217110A456BC353502D20A08",
            INIT_RAM_24 => X"28560460E9245100030C0DC251A4C1D402CC614261A2115B000411D1DA015DD0",
            INIT_RAM_25 => X"E150BB2941090150451488BC8FC501063AEC015CFC76D56C55E4A71632326293",
            INIT_RAM_26 => X"01040000259B5A62A9ACCCDE0502A0A018B190726B649948C64AD92658C1922A",
            INIT_RAM_27 => X"C848D5818383860F806126680D9037AC441004840AD4310760819046A55808E5",
            INIT_RAM_28 => X"20D183053A15555331409B059BFB6410410CC8ABD6B494944DE0A7830B150AAF",
            INIT_RAM_29 => X"123A1485B9890197750FD6AA9E0400000010000415551504545041A86AC2EB20",
            INIT_RAM_2A => X"205B3D9D0297823E748119980000820916545050BF77E6605547AECF964EE102",
            INIT_RAM_2B => X"3D007F8C502301204003B2E4508E702C2EA81209D6FABAAFA23FC2D9C95F2AE5",
            INIT_RAM_2C => X"3C6FF4EDD615D01204B26DEFD363924001E870257A3C895F91F1A3E1E55A3320",
            INIT_RAM_2D => X"AE5555B502A7F5854894C0A11594BD3E8D70C58B767050998C8DBCE48B9D1FCB",
            INIT_RAM_2E => X"E0DFC3D5EFE9CFFF43B09D340628202CE2031554847244445554D6ABEAABEBEE",
            INIT_RAM_2F => X"3D0C20468221A9E6FFEA9996ADAEC136D8824A8EDB4001A80EAAA8636C76D860",
            INIT_RAM_30 => X"CEAF2A21C40C3BCE12C191C6FFDE3D7A86600ACE99D18905A18C846FA18BAF48",
            INIT_RAM_31 => X"1CE8F7FFADFDFFEB7F376897C02D0168425BFBFFD6FEFFF48FE5908A6E533935",
            INIT_RAM_32 => X"F0A07071F12B76DF4318E73EA199B60E7ECC21D69B8AE180C8AAD020EC484611",
            INIT_RAM_33 => X"037E88EE753608120730E5543EA759DD9DB2D3715C52E9CC86A63200E5503CFA",
            INIT_RAM_34 => X"6DA7FDA97D80A29960EC0F8BE70DDA56ECA30C00706904C1348C27B28A214C02",
            INIT_RAM_35 => X"5F1F37CC47502BFDC6015E1EDDA326A6C51CF3C1F90BF3319964D3F7F3F9280F",
            INIT_RAM_36 => X"9AB36CE939D8C505D7926380E1284510EF807B2E70E3CE2DBA8577FBC238DDAB",
            INIT_RAM_37 => X"4E8A1C5554D14A124FD73F32692136B898DB3C3356D3748EE1F3EC99712C32AF",
            INIT_RAM_38 => X"C6CC08D082742C7B9C8A4186E00BAEDDA466C3924D365936D966003EC0D70698",
            INIT_RAM_39 => X"DB5BDBFED6111060952622150248737130E9AD230A82E32DAC06101D3B4B428E",
            INIT_RAM_3A => X"9EEA7DEDDD27BA52A5212180A0814001841C475661CE2084B66DB12D9B6C4B66",
            INIT_RAM_3B => X"4574449909AA2281574ABDC2AF4018098038110245A0D7EC78097700D04E83A4",
            INIT_RAM_3C => X"CCA8CEF241448805A0E251C4A504250C150615269527B51B63348F117E2C6C7C",
            INIT_RAM_3D => X"9837615FEC2937278B31E19B3B14642A1D68E50D881930D387DF99CCCC9F9E61",
            INIT_RAM_3E => X"139ACE6EBC36ACB8AD93EA23D4387D9CDD786BDA6D4ED82E049AAAAD89DCCDE5",
            INIT_RAM_3F => X"72A0000002E29E9405902E12574985A854381210B4A152970A521A861B83A528"
        )
        port map (
            DO => prom_inst_16_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_17: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"97E42BA702155AF7AB422B5B647561935CD2B6357F49C99DC983C8F6D01A728B",
            INIT_RAM_01 => X"1250010D180454827A0E040040692415D222BA8E29DCEF710B77D8FC4B52B025",
            INIT_RAM_02 => X"B653590C7D810C15C2857B460280048007FE0801004D2BA423904104201D5215",
            INIT_RAM_03 => X"0568C11050163AAA612C780C2E983DC490024315217110A456BC353502D20A08",
            INIT_RAM_04 => X"28560460E9245100030C0DC251A4C1D402CC614261A2115B000411D1DA015DD0",
            INIT_RAM_05 => X"E150BB2941090150451488BC8FC501063AEC015CFC76D56C55E4A71632326293",
            INIT_RAM_06 => X"01040000259B5A62A9ACCCDE0502A0A018B190726B649948C64AD92658C1922A",
            INIT_RAM_07 => X"C848D5818383860F806126680D9037AC441004840AD4310760819046A55808E5",
            INIT_RAM_08 => X"20D183053A15555331409B059BFB6410410CC8ABD6B494944DE0A7830B150AAF",
            INIT_RAM_09 => X"123A1485B9890197750FD6AA9E0400000010000415551504545041A86AC2EB20",
            INIT_RAM_0A => X"205B3D9D0297823E748119980000820916545050BF77E6605547AECF964EE102",
            INIT_RAM_0B => X"3D007F8C502301204003B2E4508E702C2EA81209D6FABAAFA23FC2D9C95F2AE5",
            INIT_RAM_0C => X"3C6FF4EDD615D01204B26DEFD363924001E870257A3C895F91F1A3E1E55A3320",
            INIT_RAM_0D => X"AE5555B502A7F5854894C0A11594BD3E8D70C58B767050998C8DBCE48B9D1FCB",
            INIT_RAM_0E => X"E0DFC3D5EFE9CFFF43B09D340628202CE2031554847244445554D6ABEAABEBEE",
            INIT_RAM_0F => X"3D0C20468221A9E6FFEA9996ADAEC136D8824A8EDB4001A80EAAA8636C76D860",
            INIT_RAM_10 => X"CEAF2A21C40C3BCE12C191C6FFDE3D7A86600ACE99D18905A18C846FA18BAF48",
            INIT_RAM_11 => X"1CE8F7FFADFDFFEB7F376897C02D0168425BFBFFD6FEFFF48FE5908A6E533935",
            INIT_RAM_12 => X"F0A07071F12B76DF4318E73EA199B60E7ECC21D69B8AE180C8AAD020EC484611",
            INIT_RAM_13 => X"037E88EE753608120730E5543EA759DD9DB2D3715C52E9CC86A63200E5503CFA",
            INIT_RAM_14 => X"6DA7FDA97D80A29960EC0F8BE70DDA56ECA30C00706904C1348C27B28A214C02",
            INIT_RAM_15 => X"5F1F37CC47502BFDC6015E1EDDA326A6C51CF3C1F90BF3319964D3F7F3F9280F",
            INIT_RAM_16 => X"9AB36CE939D8C505D7926380E1284510EF807B2E70E3CE2DBA8577FBC238DDAB",
            INIT_RAM_17 => X"4E8A1C5554D14A124FD73F32692136B898DB3C3356D3748EE1F3EC99712C32AF",
            INIT_RAM_18 => X"C6CC08D082742C7B9C8A4186E00BAEDDA466C3924D365936D966003EC0D70698",
            INIT_RAM_19 => X"DB5BDBFED6111060952622150248737130E9AD230A82E32DAC06101D3B4B428E",
            INIT_RAM_1A => X"9EEA7DEDDD27BA52A5212180A0814001841C475661CE2084B66DB12D9B6C4B66",
            INIT_RAM_1B => X"4574449909AA2281574ABDC2AF4018098038110245A0D7EC78097700D04E83A4",
            INIT_RAM_1C => X"CCA8CEF241448805A0E251C4A504250C150615269527B51B63348F117E2C6C7C",
            INIT_RAM_1D => X"9837615FEC2937278B31E19B3B14642A1D68E50D881930D387DF99CCCC9F9E61",
            INIT_RAM_1E => X"139ACE6EBC36ACB8AD93EA23D4387D9CDD786BDA6D4ED82E049AAAAD89DCCDE5",
            INIT_RAM_1F => X"72A0000002E29E9405902E12574985A854381210B4A152970A521A861B83A528",
            INIT_RAM_20 => X"97E42BA702155AF7AB422B5B647561935CD2B6357F49C99DC983C8F6D01A728B",
            INIT_RAM_21 => X"1250010D180454827A0E040040692415D222BA8E29DCEF710B77D8FC4B52B025",
            INIT_RAM_22 => X"B653590C7D810C15C2857B460280048007FE0801004D2BA423904104201D5215",
            INIT_RAM_23 => X"0568C11050163AAA612C780C2E983DC490024315217110A456BC353502D20A08",
            INIT_RAM_24 => X"28560460E9245100030C0DC251A4C1D402CC614261A2115B000411D1DA015DD0",
            INIT_RAM_25 => X"E150BB2941090150451488BC8FC501063AEC015CFC76D56C55E4A71632326293",
            INIT_RAM_26 => X"01040000259B5A62A9ACCCDE0502A0A018B190726B649948C64AD92658C1922A",
            INIT_RAM_27 => X"C848D5818383860F806126680D9037AC441004840AD4310760819046A55808E5",
            INIT_RAM_28 => X"20D183053A15555331409B059BFB6410410CC8ABD6B494944DE0A7830B150AAF",
            INIT_RAM_29 => X"123A1485B9890197750FD6AA9E0400000010000415551504545041A86AC2EB20",
            INIT_RAM_2A => X"205B3D9D0297823E748119980000820916545050BF77E6605547AECF964EE102",
            INIT_RAM_2B => X"3D007F8C502301204003B2E4508E702C2EA81209D6FABAAFA23FC2D9C95F2AE5",
            INIT_RAM_2C => X"3C6FF4EDD615D01204B26DEFD363924001E870257A3C895F91F1A3E1E55A3320",
            INIT_RAM_2D => X"AE5555B502A7F5854894C0A11594BD3E8D70C58B767050998C8DBCE48B9D1FCB",
            INIT_RAM_2E => X"E0DFC3D5EFE9CFFF43B09D340628202CE2031554847244445554D6ABEAABEBEE",
            INIT_RAM_2F => X"3D0C20468221A9E6FFEA9996ADAEC136D8824A8EDB4001A80EAAA8636C76D860",
            INIT_RAM_30 => X"CEAF2A21C40C3BCE12C191C6FFDE3D7A86600ACE99D18905A18C846FA18BAF48",
            INIT_RAM_31 => X"1CE8F7FFADFDFFEB7F376897C02D0168425BFBFFD6FEFFF48FE5908A6E533935",
            INIT_RAM_32 => X"F0A07071F12B76DF4318E73EA199B60E7ECC21D69B8AE180C8AAD020EC484611",
            INIT_RAM_33 => X"037E88EE753608120730E5543EA759DD9DB2D3715C52E9CC86A63200E5503CFA",
            INIT_RAM_34 => X"6DA7FDA97D80A29960EC0F8BE70DDA56ECA30C00706904C1348C27B28A214C02",
            INIT_RAM_35 => X"5F1F37CC47502BFDC6015E1EDDA326A6C51CF3C1F90BF3319964D3F7F3F9280F",
            INIT_RAM_36 => X"9AB36CE939D8C505D7926380E1284510EF807B2E70E3CE2DBA8577FBC238DDAB",
            INIT_RAM_37 => X"4E8A1C5554D14A124FD73F32692136B898DB3C3356D3748EE1F3EC99712C32AF",
            INIT_RAM_38 => X"C6CC08D082742C7B9C8A4186E00BAEDDA466C3924D365936D966003EC0D70698",
            INIT_RAM_39 => X"DB5BDBFED6111060952622150248737130E9AD230A82E32DAC06101D3B4B428E",
            INIT_RAM_3A => X"9EEA7DEDDD27BA52A5212180A0814001841C475661CE2084B66DB12D9B6C4B66",
            INIT_RAM_3B => X"4574449909AA2281574ABDC2AF4018098038110245A0D7EC78097700D04E83A4",
            INIT_RAM_3C => X"CCA8CEF241448805A0E251C4A504250C150615269527B51B63348F117E2C6C7C",
            INIT_RAM_3D => X"9837615FEC2937278B31E19B3B14642A1D68E50D881930D387DF99CCCC9F9E61",
            INIT_RAM_3E => X"139ACE6EBC36ACB8AD93EA23D4387D9CDD786BDA6D4ED82E049AAAAD89DCCDE5",
            INIT_RAM_3F => X"72A0000002E29E9405902E12574985A854381210B4A152970A521A861B83A528"
        )
        port map (
            DO => prom_inst_17_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_18: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"7697D7C6BF116E21BF42F3F0286DCF322DF7CC6360FF58848028C60002020161",
            INIT_RAM_01 => X"09C66622336C2F05B58476B69B03102ED1B10667231FD90B697E880500900934",
            INIT_RAM_02 => X"FB48C4248241AF6C248A30C41294A022E67B2280BE4C2E8C0F630E9B835ADBC9",
            INIT_RAM_03 => X"E401824DC29C331BF60FD03875500FF60CEA885D847C7E654CA839BDA0E6439A",
            INIT_RAM_04 => X"20269100004E91018481B01C01D84011104446A9224CDE0189225D310580D020",
            INIT_RAM_05 => X"565C9D63FFD367CFFEDEC4001BC652DFA84A817B40A042182188051010114808",
            INIT_RAM_06 => X"7DB5BB4C8C0641104175210B2A03C9B15989837DBA0754C5AB4FDB030A015BBE",
            INIT_RAM_07 => X"E099C4CB5A966DCC4723915A071A00413B05F58831F4723815827428BAA112E9",
            INIT_RAM_08 => X"124E7D1665A78E954E894BEF0DA3F9375CED5AAD799EC3F13589086846A1DCEE",
            INIT_RAM_09 => X"8DD2200D8DB74EFE6666776CF4E8E9B81C780C0234465A78C18DB87AC3C41964",
            INIT_RAM_0A => X"C30A1FF622806700BF282A8FC521141906C24E8DF6C429FFD7E0AAD5B0402769",
            INIT_RAM_0B => X"8E1FCE1FFAD5877D6B0586C600DAC90614011114A3602B6918D1FF24C1202968",
            INIT_RAM_0C => X"53D28DEF45AA8E0368F96596DF44CDA36C61B2681584016F7D680484EDCE0BB5",
            INIT_RAM_0D => X"00900044444044B0422017EC0540503069B55109BD085B40C20D52A86B568320",
            INIT_RAM_0E => X"1B1C72516E66266A118190AA9569585AC2B42B51A82DE6ADAB5259A67F0B0280",
            INIT_RAM_0F => X"BE856D4A0844790C6F08C9357C8E3D810491189CAB128320282A2828282B6C51",
            INIT_RAM_10 => X"1044514155410140441055005171189CAB1C844045B6075657A0847AB440C4CA",
            INIT_RAM_11 => X"689322B6018AB6DD5856F4E231C76800E39EC000005555554000554015054145",
            INIT_RAM_12 => X"425ACB9B7032518D87C7A18FB415D55864F790FA12147B13A9C4E27BC194CE94",
            INIT_RAM_13 => X"0603E32BF4681D1301A9A91C1742A988F67621C7878C6D91B88CAEDE18D000C7",
            INIT_RAM_14 => X"C6DE919F38298DE6F486671C667033C56C59C67CE448E4B39CA705F1234CF9C1",
            INIT_RAM_15 => X"336663900FB20A884180C008902114D44B0F46C7C69E9A6F0701010FAAEE8DDE",
            INIT_RAM_16 => X"3CE87FFCD4F4F7A2BDBF10610BA80C8BB1981862A804E0D4C1AC286083D39677",
            INIT_RAM_17 => X"C8CC3261B10E27BC7EB4A92602308980020641249882691A088288293210B431",
            INIT_RAM_18 => X"8C80DB032380C8E0991A731304C7B79955510E4A290ACEF926A926146C8194D9",
            INIT_RAM_19 => X"9D144A0F8F6EE0311ED271A1249939032C9F294DD9FF4B641D244F8065011889",
            INIT_RAM_1A => X"6D309835E34A14C009C0A522C4E4904E389E229E221BC78F43336E08D4C3CC11",
            INIT_RAM_1B => X"7A8C194A8E99A618F66F49331804D69411AA03B04664E84E8123B0761B410E98",
            INIT_RAM_1C => X"4552218B6DDF7DAC25A6E2B10333868036FBC1054763D2A386DE951DEA6CA545",
            INIT_RAM_1D => X"FF1C5D24349E464423A1336D9ED6DC45696FDB452C51EFBEC0CB1911D0C43562",
            INIT_RAM_1E => X"7DD0518FFCAFB07F1C4798FF1D993DB1E490D26E4532230909F0FF148FF19D93",
            INIT_RAM_1F => X"DFF7D7BE593AEF953259FF5445696D64B25CC9031CF6A6C7B0EEA6EA71FF95F4",
            INIT_RAM_20 => X"34862D1420452E49614AB6A7FF8B7DADBC5AC9F6EC92DE4C58F981B0F984DF7B",
            INIT_RAM_21 => X"660281450A4520A0C244D504062224C209523A8138449A91851FF801A021F4A4",
            INIT_RAM_22 => X"98206BAA288AA81E0ED2A365CC198C80C7092D19B826CC8061444B4A8048C942",
            INIT_RAM_23 => X"92E05F7A6108427EA301C04A8367A015A80003CC14654090498405E12235DDA4",
            INIT_RAM_24 => X"4AD53E08D847808D887F9BB4E5B0514202151AA6BE8CAF7777776C45F657EECF",
            INIT_RAM_25 => X"C089A84691934A84011411933680B82490043F7C2400080092BE2127B0829629",
            INIT_RAM_26 => X"34A15BA93D1415042214130C4AD000A292214088FD3850001534800046B82668",
            INIT_RAM_27 => X"00154AA90A3102A62C491E8C41205A523A408F0160E50046F620D4752032200C",
            INIT_RAM_28 => X"5231AAD500C0360C8542C2A24058A009480862191019A02C226CA6C509B4309B",
            INIT_RAM_29 => X"2A820680AC0599A992004ACCD4D2004AAD60430461840685A74202D082771631",
            INIT_RAM_2A => X"6AAA1682682D22E0EB0A85707185682B0150AE505E2C3A479515AB063158424B",
            INIT_RAM_2B => X"4A95A40C8191D1D4794235444063501ABD1D5C752A69876C040C4E87C20CD2D5",
            INIT_RAM_2C => X"DDA42144E85EC11980F6DA42304652331DA3314A74519D0E0233DF14854AD3A9",
            INIT_RAM_2D => X"28128819B10A00A32063807C04A3000F6A8C002001076A164AA083B251C12019",
            INIT_RAM_2E => X"00001E31B0138961ED074F6D8DA33A10C2C635C3E2CB0D719A80D9A312C7C8F8",
            INIT_RAM_2F => X"932241595832525649B322C58FA65A182B1828501AC032028F310DA124300000",
            INIT_RAM_30 => X"F0CED96D6FB0635793A1448308CD200C95514A09064B411932150C9A92290483",
            INIT_RAM_31 => X"18D90194183705B1BDE595200029E34829019E447A60768C398DAA988EF90781",
            INIT_RAM_32 => X"8B5C98298FFFFFFD1B1341A7E86DB26AEA4988AA9832EC0CCD96D6FB0E7B2287",
            INIT_RAM_33 => X"2BD6CDF633A77EAE8496855E1C6A7DF5FBD4AE98783839610FB2AE72DDBF7323",
            INIT_RAM_34 => X"B10D012B52D439CE9F08B4CDDBC8B096B77DF7DC4CACAE867A7C6CFC218466DE",
            INIT_RAM_35 => X"305C56125127C31AE04080C49736E807DED9C6E8AE4C01CDE9405F896E39D1F3",
            INIT_RAM_36 => X"1C0A30EEEAD105B466846C638AEA4A4600405EAD558AAB15291222D1222C1225",
            INIT_RAM_37 => X"A6AA95AA9EC1958BFE59FE0624240C4004E82C8F0191C4399F6BF8A80A8D8D1B",
            INIT_RAM_38 => X"2CC0A7A65892495C1DA31B5AF934E4DD24B269A92029482CDB66978A49243FC2",
            INIT_RAM_39 => X"F4A7562101474D447CB986961B1C0BE7F4D3606406137666318B33A985032139",
            INIT_RAM_3A => X"3E3103522234D59C2E0DB0F06B9FAE6481010E9C65C76534D4C2D04D8357B684",
            INIT_RAM_3B => X"3E307CBFF4C35186A524AAAC1F574368043404CF998EFC9D110E043D8C106100",
            INIT_RAM_3C => X"9197AB44EC6A8DEEAC88D68984D59A6D59320AAA6F5BFF4E0A85568CF1414162",
            INIT_RAM_3D => X"9FD9FD8596FECBC923889E2E5B6A8DC18E8BC66C1BB66DC76EA9CCFB1CCC8DED",
            INIT_RAM_3E => X"236B5B6BCDB68556AEAB0C47B6E40D769516A1173A9FCFA6A7ABB50CF6DB96D1",
            INIT_RAM_3F => X"02081AC47C549FFB71D4D4F4FCDCFB7B077305153C9190FF959B721122EF8B52"
        )
        port map (
            DO => prom_inst_18_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_2,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_19: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"111F830F9851184101370588A06D3BF9AE621E7FCE63326799C8FEFAAEFE769D",
            INIT_RAM_01 => X"EC2A08157331C6CC0E30884244916A0DE26D4D22454091290404A492016887E2",
            INIT_RAM_02 => X"96968460CA3388A03ECB45F2C4B70F1829221000FFFC7FEC346F079F13079798",
            INIT_RAM_03 => X"2251A60725008AAA056591C4000BB48C0BC29B8034A03400027B84769B520D91",
            INIT_RAM_04 => X"C13E7C640F364509212AE9CC14296E30DEA3057B35C641762CD00D40DABC2747",
            INIT_RAM_05 => X"861F8BC1993560946D92D1C0C7F046A245B5849CB751FF15B97FCD50BC7B8524",
            INIT_RAM_06 => X"E90C8E38C8E0478AD8B388F94891C9673A50BC32478E083074657E8E0EA53BEE",
            INIT_RAM_07 => X"17A24D2C636ED2478B5AE1C99D40761B1E7AA6A89DDD1BBD8DBD223E70531BCD",
            INIT_RAM_08 => X"470542C2E3C783A4C24767084C52DC209D60E95DBC096D9A0171A12D5AB99BAB",
            INIT_RAM_09 => X"5686C6CA41B2224C88D8456C1DBF20DC20A6649774CB11B69933246E9739C998",
            INIT_RAM_0A => X"3488480610A91A851E84FF08783F81AEA52D2FDC2200BC2FE81C0357FBEC1D87",
            INIT_RAM_0B => X"1620D1A60A901095D12A0973B95E20838001330138991361967847D42901910A",
            INIT_RAM_0C => X"8A370D60A0AA3E7288F4B0869FA5E703D1AE17C0EC276B2AFB747B550A8B4102",
            INIT_RAM_0D => X"95D23A0E191EBC2134B833D53D37E42B05018289A10300A188E315CE98640F54",
            INIT_RAM_0E => X"DCB42E8E77212A58842051A078007109A0D820166B8810426002844031430482",
            INIT_RAM_0F => X"C82B30679933680037A65978674DDEC2D30EEEDA78F5F2A1DEE660FFEA11B175",
            INIT_RAM_10 => X"C194E3598360AFB031A1690F4625BB628363B4C90A400E3A04DAA70DA0CC3776",
            INIT_RAM_11 => X"9DD952B29003D7767BA581A68BC41C2B16AD6EB57F1D048CD4E464190D25ADF2",
            INIT_RAM_12 => X"3B9AF0147BDB7730B4E11D9D11C1D0C3C6E0B6F242719988ACDDB17B4D81882E",
            INIT_RAM_13 => X"C653A0510A1B00C36AC88058CAC126E14E198DFB07E80C3EC1510BB08F8F851C",
            INIT_RAM_14 => X"1310B00A49902C0104004C654E0582040001103654011012021912281216B000",
            INIT_RAM_15 => X"A2E5A64B241400267194CD524499BC01D31058CD18684A817A5800B65143281C",
            INIT_RAM_16 => X"A0CC44CC94E2649242CE08191634113154562B149100204551178DE805D98EC8",
            INIT_RAM_17 => X"1AA1C248D293110CB951445117D9B6AA500F65068B8CC508BD00184F8501B010",
            INIT_RAM_18 => X"89B6054CC727D292805705A932685B6A31111371390B240EC3CC85D331813EB1",
            INIT_RAM_19 => X"316412C4900F646A36630261DA093053D98F19D2C5B653195D4A71AA5682B29B",
            INIT_RAM_1A => X"08980020680249882691A6C0488292310B4313CE87FFCD5329A64B708CAC8533",
            INIT_RAM_1B => X"2760A263DBCCAAA88712242B3BE49AA4938990229B391158C726BC7EB4ECC323",
            INIT_RAM_1C => X"F10410AC463BF80C9074917E0674A12830EFA280EBD3131E484A255D0191C685",
            INIT_RAM_1D => X"3DA2C64840C2CCE811522B42008095E5A456C98F4B25EAEA410610545024640C",
            INIT_RAM_1E => X"7888672DC999B7046A61E60810A7434450E3D33E330F321A18E8A120D1EDC862",
            INIT_RAM_1F => X"35861A00A6112A1481AF1A50A6004A05291627227FF08229B87389E08119A28A",
            INIT_RAM_20 => X"4B710C9DC948F06010DF01D880C4444BE8854062D10DD93F30A62AA7FD227C4C",
            INIT_RAM_21 => X"5BFE5CE861A20F71E8032916A78F29CC546518461522E4E14998DD54BC0E40B6",
            INIT_RAM_22 => X"40B6C18000680080125C75401AEC44E8C01A8D40D1412B25A09F7600B0C6FEC6",
            INIT_RAM_23 => X"7000000030082004A17800828F090A0C318CE120012172286317922341A2A128",
            INIT_RAM_24 => X"093E11673256B3169C12284980E92A034141E0782507800F8100009C403C0786",
            INIT_RAM_25 => X"8249144AB52CED94200A0202A88510084D938A30A34512C0CE098F08A98900F2",
            INIT_RAM_26 => X"AB6AA38578BD55CEC9AA28082C285B8C0201104838AD512AC160C13C70620B81",
            INIT_RAM_27 => X"1228D91C352915424000000AA0088F63153A8AD81B945C8789F01C86548D12CE",
            INIT_RAM_28 => X"9A22242CB58413089465B246231330D806105010035100B08761A08506094160",
            INIT_RAM_29 => X"00CC60799124A8520C08050122171281808058018C38A645D07931896B39ED25",
            INIT_RAM_2A => X"3C251301FB2CA45562245308885131119115C652B2493252340201101942D260",
            INIT_RAM_2B => X"2A086B442661015380041594608092D9CB919250100A37DDA3919A1427F66096",
            INIT_RAM_2C => X"02288A804612A2A0A102A418CBDFBA554499541660F812464011010126314289",
            INIT_RAM_2D => X"6059E332C311521E6522901852D484B423A98816C9B26A08C92368E9F8055245",
            INIT_RAM_2E => X"35188757AC5A42DEB501FE010586249AC1EA60D08F4267D2843763CFC9190C05",
            INIT_RAM_2F => X"E2975A2686A7AE0288F140141B698E2A82A835F478453A1D722CFCED12859FD7",
            INIT_RAM_30 => X"8DC6A06905054C8C36E4199E74638E6532965218A965909BA456000451343351",
            INIT_RAM_31 => X"7BB16DDB96B7845371C30B55DB96C8F6EB4B453242FF6A4DF84A76B5AEDC88A6",
            INIT_RAM_32 => X"FF7FFF7D5712524D4A30723514B2B3064A84B4742D484152FB611117AA9D9B7E",
            INIT_RAM_33 => X"0E78522BA2812C1454A502ED1A59CBD76A034756F5765DF7555F57575F7F57FF",
            INIT_RAM_34 => X"F88D5002628FFD13203066C850F10649F21319109208387641120B362124803F",
            INIT_RAM_35 => X"52979565817114DE46462844A57F7958873FC4B255C8AE549BDD1A87415D5018",
            INIT_RAM_36 => X"453FDC2219C225E421B320085A8FBFD0C42135B16448DFC226E09B3438A740C3",
            INIT_RAM_37 => X"5861917919344A4685CC0990862A11324792E761B6D41C0FCC0838C1C27211A2",
            INIT_RAM_38 => X"B28480C32660C60C6D1A6AA9048E925F15015010D2195982823226DED0ADFCB8",
            INIT_RAM_39 => X"B88334AA071AA818B16C242E6496AD88425096D575AD8A1A2E7A8971313EE1B1",
            INIT_RAM_3A => X"9BB9F1C12F200009D3425B5486BE6A5A1183286713CA207720DD42E52C8FC903",
            INIT_RAM_3B => X"8000000125CC06AF3BB0A68881710C814B500D182A48301C0FC0001EE0E1E5C7",
            INIT_RAM_3C => X"000000000000000000000000006EF6B03EB643C2A5704C696AB9AFD1DFFFDB69",
            INIT_RAM_3D => X"024428106448524A624A4A24425242522060108010543C00044A105424005E00",
            INIT_RAM_3E => X"807E7E10005270182040407E4A1252124208084008404208420A4A42424A125A",
            INIT_RAM_3F => X"A50276000854A0103840403E540424244404783E18807A08A47C54484448544A"
        )
        port map (
            DO => prom_inst_19_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_20: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"1EA06DB51F7E00FFE0037F017B861FE79F7CFF16FC9828104EC4DF8940580883",
            INIT_RAM_01 => X"5B50294907F75E7BAD74549269BA592524BBDD5ECFDEFFD4B3D2752DED50F05D",
            INIT_RAM_02 => X"24579159100A40B9908EDB8C0A50C0443C5A2B30CC4108A4DD404C0445CC4225",
            INIT_RAM_03 => X"C55ACB2C902EDFE85CD96209973E6DADFA174BB937EB7AB4F9EB8C4C19A85021",
            INIT_RAM_04 => X"0A578EA3320F6A4001188B66679E9E822FE80A51883A9EDA029E87ED6526A3E5",
            INIT_RAM_05 => X"8B922D5E48A414150104001298800A413429DD98B4EDD5F565DCDA69AEBDA6D7",
            INIT_RAM_06 => X"0B9EE0FE00000007FB2EEEDEAA1FFFF1734D75FDAD6B78B6A7B35ADE26B9EC4C",
            INIT_RAM_07 => X"110AD5059683765A82E7EAEA2D5EB6FA4A9284865E50E9355D9498E7FE156A82",
            INIT_RAM_08 => X"04C3815132A10410C4133901BBB7E000821219387E698B8849600063EF5D9FAC",
            INIT_RAM_09 => X"5AF036B7AB7D8FBBAE17AF65FF515555555555440000E8A5001501084238DB20",
            INIT_RAM_0A => X"C113D231DE3E262F6F2133354C14BEFD94E05882526BEF915EB9ADDFC44CFF2B",
            INIT_RAM_0B => X"FD8F11F4DBF6A43160FCEFEC54EC6BCF5D30FB1B07F5CDEF8AF2164983605B40",
            INIT_RAM_0C => X"DF5FFBF5AFEBA087FBFC0ABF47AAF515358D565BFBD8CAD467F28E7963570482",
            INIT_RAM_0D => X"570165302B27F9C963A579352088DE292816FA24A588D0AAAA825CAA32D46EEB",
            INIT_RAM_0E => X"B033ABFBF6D7D6DB774D5ABDFFF502AED6531FF8847B5543C446D7BBFA2ABAAC",
            INIT_RAM_0F => X"BDFFBBFF502BF566FF809BADDB6A407FF82E8027FF7FFE700C888BDFF13FFFDA",
            INIT_RAM_10 => X"99EE454406AABE080381818FFF5EADFFBC2C00AFFD2780DC7D0B000D83FA1F75",
            INIT_RAM_11 => X"548EF7FFADB5FFEB6D5B6ADA51D050DD7F000124800049214AA6A25F7E2A663D",
            INIT_RAM_12 => X"F156800D700A00090739CE7809B9DA1D5A0092810760D3AD1DDEDABAFA240101",
            INIT_RAM_13 => X"8762FB9177347FFA5E108004AC101329E81020EC1A508009101EBBB5000408FE",
            INIT_RAM_14 => X"009249296016F2779291A9ABC031415E222FBF57C42B5710A9B85DFE9E1CC537",
            INIT_RAM_15 => X"C470FC3BDFBEAC5D5DE900E24417D2D85571ACE0F47D7A9B394201248292A5BE",
            INIT_RAM_16 => X"9DB404D421B08FFF0040224C08ABEA952F005D45135346F95DE551B98EE145F4",
            INIT_RAM_17 => X"6D5450F7FE83F71468137408048326BD04920D523697404D07820049356A36AA",
            INIT_RAM_18 => X"020BD927016E78FA948D8928017A8124124E821D80020009018155051AFF5200",
            INIT_RAM_19 => X"92000124800807652B490357B084A40404006452A2C7AC64A245E9B05003AA80",
            INIT_RAM_1A => X"6F5249868A5BD4601989D92E84DD3CA4A6566548939CE7000049200012480004",
            INIT_RAM_1B => X"CB77CC9DB37F75C86ADCDE37379FEE102044FFBFE370E7DE42B1A2D8E0399767",
            INIT_RAM_1C => X"80AF451F7BCD9A2F65F673E8A5983D9E7D96BD82AD3BA97B0A9C8B99BE08CC58",
            INIT_RAM_1D => X"C054016F8408AB11E00B035BA113584C0568DBF6EFF552D6031C9E4D001F5EE9",
            INIT_RAM_1E => X"2302A45530B532E1AA258F417C7ABD48AA616DEB4E4CC016451CCCCE48011127",
            INIT_RAM_1F => X"5A900000055B6F2605B7FF21DF8A070204001039C003A7B8257D58201B62C8BD",
            INIT_RAM_20 => X"1EA06DB51F7E00FFE0037F017B861FE79F7CFF16FC9828104EC4DF8940580883",
            INIT_RAM_21 => X"5B50294907F75E7BAD74549269BA592524BBDD5ECFDEFFD4B3D2752DED50F05D",
            INIT_RAM_22 => X"24579159100A40B9908EDB8C0A50C0443C5A2B30CC4108A4DD404C0445CC4225",
            INIT_RAM_23 => X"C55ACB2C902EDFE85CD96209973E6DADFA174BB937EB7AB4F9EB8C4C19A85021",
            INIT_RAM_24 => X"0A578EA3320F6A4001188B66679E9E822FE80A51883A9EDA029E87ED6526A3E5",
            INIT_RAM_25 => X"8B922D5E48A414150104001298800A413429DD98B4EDD5F565DCDA69AEBDA6D7",
            INIT_RAM_26 => X"0B9EE0FE00000007FB2EEEDEAA1FFFF1734D75FDAD6B78B6A7B35ADE26B9EC4C",
            INIT_RAM_27 => X"110AD5059683765A82E7EAEA2D5EB6FA4A9284865E50E9355D9498E7FE156A82",
            INIT_RAM_28 => X"04C3815132A10410C4133901BBB7E000821219387E698B8849600063EF5D9FAC",
            INIT_RAM_29 => X"5AF036B7AB7D8FBBAE17AF65FF515555555555440000E8A5001501084238DB20",
            INIT_RAM_2A => X"C113D231DE3E262F6F2133354C14BEFD94E05882526BEF915EB9ADDFC44CFF2B",
            INIT_RAM_2B => X"FD8F11F4DBF6A43160FCEFEC54EC6BCF5D30FB1B07F5CDEF8AF2164983605B40",
            INIT_RAM_2C => X"DF5FFBF5AFEBA087FBFC0ABF47AAF515358D565BFBD8CAD467F28E7963570482",
            INIT_RAM_2D => X"570165302B27F9C963A579352088DE292816FA24A588D0AAAA825CAA32D46EEB",
            INIT_RAM_2E => X"B033ABFBF6D7D6DB774D5ABDFFF502AED6531FF8847B5543C446D7BBFA2ABAAC",
            INIT_RAM_2F => X"BDFFBBFF502BF566FF809BADDB6A407FF82E8027FF7FFE700C888BDFF13FFFDA",
            INIT_RAM_30 => X"99EE454406AABE080381818FFF5EADFFBC2C00AFFD2780DC7D0B000D83FA1F75",
            INIT_RAM_31 => X"548EF7FFADB5FFEB6D5B6ADA51D050DD7F000124800049214AA6A25F7E2A663D",
            INIT_RAM_32 => X"F156800D700A00090739CE7809B9DA1D5A0092810760D3AD1DDEDABAFA240101",
            INIT_RAM_33 => X"8762FB9177347FFA5E108004AC101329E81020EC1A508009101EBBB5000408FE",
            INIT_RAM_34 => X"009249296016F2779291A9ABC031415E222FBF57C42B5710A9B85DFE9E1CC537",
            INIT_RAM_35 => X"C470FC3BDFBEAC5D5DE900E24417D2D85571ACE0F47D7A9B394201248292A5BE",
            INIT_RAM_36 => X"9DB404D421B08FFF0040224C08ABEA952F005D45135346F95DE551B98EE145F4",
            INIT_RAM_37 => X"6D5450F7FE83F71468137408048326BD04920D523697404D07820049356A36AA",
            INIT_RAM_38 => X"020BD927016E78FA948D8928017A8124124E821D80020009018155051AFF5200",
            INIT_RAM_39 => X"92000124800807652B490357B084A40404006452A2C7AC64A245E9B05003AA80",
            INIT_RAM_3A => X"6F5249868A5BD4601989D92E84DD3CA4A6566548939CE7000049200012480004",
            INIT_RAM_3B => X"CB77CC9DB37F75C86ADCDE37379FEE102044FFBFE370E7DE42B1A2D8E0399767",
            INIT_RAM_3C => X"80AF451F7BCD9A2F65F673E8A5983D9E7D96BD82AD3BA97B0A9C8B99BE08CC58",
            INIT_RAM_3D => X"C054016F8408AB11E00B035BA113584C0568DBF6EFF552D6031C9E4D001F5EE9",
            INIT_RAM_3E => X"2302A45530B532E1AA258F417C7ABD48AA616DEB4E4CC016451CCCCE48011127",
            INIT_RAM_3F => X"5A900000055B6F2605B7FF21DF8A070204001039C003A7B8257D58201B62C8BD"
        )
        port map (
            DO => prom_inst_20_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_21: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"1EA06DB51F7E00FFE0037F017B861FE79F7CFF16FC9828104EC4DF8940580883",
            INIT_RAM_01 => X"5B50294907F75E7BAD74549269BA592524BBDD5ECFDEFFD4B3D2752DED50F05D",
            INIT_RAM_02 => X"24579159100A40B9908EDB8C0A50C0443C5A2B30CC4108A4DD404C0445CC4225",
            INIT_RAM_03 => X"C55ACB2C902EDFE85CD96209973E6DADFA174BB937EB7AB4F9EB8C4C19A85021",
            INIT_RAM_04 => X"0A578EA3320F6A4001188B66679E9E822FE80A51883A9EDA029E87ED6526A3E5",
            INIT_RAM_05 => X"8B922D5E48A414150104001298800A413429DD98B4EDD5F565DCDA69AEBDA6D7",
            INIT_RAM_06 => X"0B9EE0FE00000007FB2EEEDEAA1FFFF1734D75FDAD6B78B6A7B35ADE26B9EC4C",
            INIT_RAM_07 => X"110AD5059683765A82E7EAEA2D5EB6FA4A9284865E50E9355D9498E7FE156A82",
            INIT_RAM_08 => X"04C3815132A10410C4133901BBB7E000821219387E698B8849600063EF5D9FAC",
            INIT_RAM_09 => X"5AF036B7AB7D8FBBAE17AF65FF515555555555440000E8A5001501084238DB20",
            INIT_RAM_0A => X"C113D231DE3E262F6F2133354C14BEFD94E05882526BEF915EB9ADDFC44CFF2B",
            INIT_RAM_0B => X"FD8F11F4DBF6A43160FCEFEC54EC6BCF5D30FB1B07F5CDEF8AF2164983605B40",
            INIT_RAM_0C => X"DF5FFBF5AFEBA087FBFC0ABF47AAF515358D565BFBD8CAD467F28E7963570482",
            INIT_RAM_0D => X"570165302B27F9C963A579352088DE292816FA24A588D0AAAA825CAA32D46EEB",
            INIT_RAM_0E => X"B033ABFBF6D7D6DB774D5ABDFFF502AED6531FF8847B5543C446D7BBFA2ABAAC",
            INIT_RAM_0F => X"BDFFBBFF502BF566FF809BADDB6A407FF82E8027FF7FFE700C888BDFF13FFFDA",
            INIT_RAM_10 => X"99EE454406AABE080381818FFF5EADFFBC2C00AFFD2780DC7D0B000D83FA1F75",
            INIT_RAM_11 => X"548EF7FFADB5FFEB6D5B6ADA51D050DD7F000124800049214AA6A25F7E2A663D",
            INIT_RAM_12 => X"F156800D700A00090739CE7809B9DA1D5A0092810760D3AD1DDEDABAFA240101",
            INIT_RAM_13 => X"8762FB9177347FFA5E108004AC101329E81020EC1A508009101EBBB5000408FE",
            INIT_RAM_14 => X"009249296016F2779291A9ABC031415E222FBF57C42B5710A9B85DFE9E1CC537",
            INIT_RAM_15 => X"C470FC3BDFBEAC5D5DE900E24417D2D85571ACE0F47D7A9B394201248292A5BE",
            INIT_RAM_16 => X"9DB404D421B08FFF0040224C08ABEA952F005D45135346F95DE551B98EE145F4",
            INIT_RAM_17 => X"6D5450F7FE83F71468137408048326BD04920D523697404D07820049356A36AA",
            INIT_RAM_18 => X"020BD927016E78FA948D8928017A8124124E821D80020009018155051AFF5200",
            INIT_RAM_19 => X"92000124800807652B490357B084A40404006452A2C7AC64A245E9B05003AA80",
            INIT_RAM_1A => X"6F5249868A5BD4601989D92E84DD3CA4A6566548939CE7000049200012480004",
            INIT_RAM_1B => X"CB77CC9DB37F75C86ADCDE37379FEE102044FFBFE370E7DE42B1A2D8E0399767",
            INIT_RAM_1C => X"80AF451F7BCD9A2F65F673E8A5983D9E7D96BD82AD3BA97B0A9C8B99BE08CC58",
            INIT_RAM_1D => X"C054016F8408AB11E00B035BA113584C0568DBF6EFF552D6031C9E4D001F5EE9",
            INIT_RAM_1E => X"2302A45530B532E1AA258F417C7ABD48AA616DEB4E4CC016451CCCCE48011127",
            INIT_RAM_1F => X"5A900000055B6F2605B7FF21DF8A070204001039C003A7B8257D58201B62C8BD",
            INIT_RAM_20 => X"1EA06DB51F7E00FFE0037F017B861FE79F7CFF16FC9828104EC4DF8940580883",
            INIT_RAM_21 => X"5B50294907F75E7BAD74549269BA592524BBDD5ECFDEFFD4B3D2752DED50F05D",
            INIT_RAM_22 => X"24579159100A40B9908EDB8C0A50C0443C5A2B30CC4108A4DD404C0445CC4225",
            INIT_RAM_23 => X"C55ACB2C902EDFE85CD96209973E6DADFA174BB937EB7AB4F9EB8C4C19A85021",
            INIT_RAM_24 => X"0A578EA3320F6A4001188B66679E9E822FE80A51883A9EDA029E87ED6526A3E5",
            INIT_RAM_25 => X"8B922D5E48A414150104001298800A413429DD98B4EDD5F565DCDA69AEBDA6D7",
            INIT_RAM_26 => X"0B9EE0FE00000007FB2EEEDEAA1FFFF1734D75FDAD6B78B6A7B35ADE26B9EC4C",
            INIT_RAM_27 => X"110AD5059683765A82E7EAEA2D5EB6FA4A9284865E50E9355D9498E7FE156A82",
            INIT_RAM_28 => X"04C3815132A10410C4133901BBB7E000821219387E698B8849600063EF5D9FAC",
            INIT_RAM_29 => X"5AF036B7AB7D8FBBAE17AF65FF515555555555440000E8A5001501084238DB20",
            INIT_RAM_2A => X"C113D231DE3E262F6F2133354C14BEFD94E05882526BEF915EB9ADDFC44CFF2B",
            INIT_RAM_2B => X"FD8F11F4DBF6A43160FCEFEC54EC6BCF5D30FB1B07F5CDEF8AF2164983605B40",
            INIT_RAM_2C => X"DF5FFBF5AFEBA087FBFC0ABF47AAF515358D565BFBD8CAD467F28E7963570482",
            INIT_RAM_2D => X"570165302B27F9C963A579352088DE292816FA24A588D0AAAA825CAA32D46EEB",
            INIT_RAM_2E => X"B033ABFBF6D7D6DB774D5ABDFFF502AED6531FF8847B5543C446D7BBFA2ABAAC",
            INIT_RAM_2F => X"BDFFBBFF502BF566FF809BADDB6A407FF82E8027FF7FFE700C888BDFF13FFFDA",
            INIT_RAM_30 => X"99EE454406AABE080381818FFF5EADFFBC2C00AFFD2780DC7D0B000D83FA1F75",
            INIT_RAM_31 => X"548EF7FFADB5FFEB6D5B6ADA51D050DD7F000124800049214AA6A25F7E2A663D",
            INIT_RAM_32 => X"F156800D700A00090739CE7809B9DA1D5A0092810760D3AD1DDEDABAFA240101",
            INIT_RAM_33 => X"8762FB9177347FFA5E108004AC101329E81020EC1A508009101EBBB5000408FE",
            INIT_RAM_34 => X"009249296016F2779291A9ABC031415E222FBF57C42B5710A9B85DFE9E1CC537",
            INIT_RAM_35 => X"C470FC3BDFBEAC5D5DE900E24417D2D85571ACE0F47D7A9B394201248292A5BE",
            INIT_RAM_36 => X"9DB404D421B08FFF0040224C08ABEA952F005D45135346F95DE551B98EE145F4",
            INIT_RAM_37 => X"6D5450F7FE83F71468137408048326BD04920D523697404D07820049356A36AA",
            INIT_RAM_38 => X"020BD927016E78FA948D8928017A8124124E821D80020009018155051AFF5200",
            INIT_RAM_39 => X"92000124800807652B490357B084A40404006452A2C7AC64A245E9B05003AA80",
            INIT_RAM_3A => X"6F5249868A5BD4601989D92E84DD3CA4A6566548939CE7000049200012480004",
            INIT_RAM_3B => X"CB77CC9DB37F75C86ADCDE37379FEE102044FFBFE370E7DE42B1A2D8E0399767",
            INIT_RAM_3C => X"80AF451F7BCD9A2F65F673E8A5983D9E7D96BD82AD3BA97B0A9C8B99BE08CC58",
            INIT_RAM_3D => X"C054016F8408AB11E00B035BA113584C0568DBF6EFF552D6031C9E4D001F5EE9",
            INIT_RAM_3E => X"2302A45530B532E1AA258F417C7ABD48AA616DEB4E4CC016451CCCCE48011127",
            INIT_RAM_3F => X"5A900000055B6F2605B7FF21DF8A070204001039C003A7B8257D58201B62C8BD"
        )
        port map (
            DO => prom_inst_21_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_22: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"5ED5446F7F03EA49CF4B3E70847C734C2E69C89C94F3F917330F3F03010101ED",
            INIT_RAM_01 => X"ED3499F805925BEB6E4E5DDBAD45EEB3E925E4445C965C31ED54A90082490012",
            INIT_RAM_02 => X"51A8ED44B6712D9265512A8DB7BDE90B797B1C52DC172E956F63805B2E6C93B6",
            INIT_RAM_03 => X"C080C18DE6283556C90B22548121816D80AACBD649FCED00104732EE8B79D392",
            INIT_RAM_04 => X"FFF7FFFEFFEFFFFDFFFEFC3FFF7E0414150507FA7D832182530C3CDAFB772A45",
            INIT_RAM_05 => X"EBA71048B2C4972B37E7D00005004AC0DBFDFEFFFFFFBFFBFFFDFFF7FFFBFFFD",
            INIT_RAM_06 => X"54A4450EBB205541150ADD6FD3A754352A592C72154FEC92128A64CCAD258547",
            INIT_RAM_07 => X"E38D332F1AAEDDEB050293FC07321EFBBFAE37D8D9B452283FC0737DEF0BBBFD",
            INIT_RAM_08 => X"407B451F34F1BE9EC1DC6AAC196B896C5548D2690AAC06B470554A5D55A9BBBE",
            INIT_RAM_09 => X"01F4F0092925E45444C45544BBAC8D3008CCEB272544CA7208D92A2B6B606BB0",
            INIT_RAM_0A => X"D83C79BEAE8244530040221D8049D0950FFFD11FBFDC00B2D7A622851872EEE5",
            INIT_RAM_0B => X"249A240D26AD27095A41268494189A1028612050A6C14242D586EF0929304A18",
            INIT_RAM_0C => X"02CA082704201E606081041083042187FFC64BB97FFDE1431C608300A96A82AD",
            INIT_RAM_0D => X"00D80050504505E400F1637EF1E21260C9E1D68507C42B035208FAE8284606A4",
            INIT_RAM_0E => X"7955548A4B7F493C9D0950888141F839C271084852092129215ED124762C0409",
            INIT_RAM_0F => X"A3BBB6B4801D051EFC4E8B4A8A8CF7AB5FC4D4802A4A16A2A2A0A2A2A2A04A95",
            INIT_RAM_10 => X"0541451044514155410100445044D4802A4A840277FE96BE1C4801CDF0CB0402",
            INIT_RAM_11 => X"264C9B1E068C1E788863F6E929274554924E8000000000001555554000554015",
            INIT_RAM_12 => X"9017643DA8D558A45B6EC95D5933173255B3584D4F0B9A56D269349A64A35873",
            INIT_RAM_13 => X"0E4DA3FA8C8E6C3269D578C52F0BE920E9A9199B5B2592AE4465F7360B2C55FB",
            INIT_RAM_14 => X"2491462C24A169148A318B7118B6C2DC4891285B8ABEACAAD664137325F0B77E",
            INIT_RAM_15 => X"065357299DA40BF4AAE5E99E3A93A9AA149E0AC5ECBCD65DAE4399B607492931",
            INIT_RAM_16 => X"328F4006D2EDA14C3FD4A275A7AD1D3732CC1D4BAD0D4E8EC9144EFBA3C59E71",
            INIT_RAM_17 => X"6020EDD89AFD20B71CDCC482411210806202DB0249080008652640248108806A",
            INIT_RAM_18 => X"421F25E9D24A749004207A124906B066A8A1A94A9B34B886CF62A4908840DC4F",
            INIT_RAM_19 => X"FABEC93A5C919926792E545DB6D6842A176CD90554E6D737D24AF39464484E64",
            INIT_RAM_1A => X"16BA417F77BD7723BE2FFF2F6CA5928C9FBD086787B0F5D292DA89B72257210C",
            INIT_RAM_1B => X"332A6323484AD309FA866688C0DDCBC979A3D2B8A0083C83CCCDC2C905A58164",
            INIT_RAM_1C => X"C108B64A4A9249061A1AFF1AA4261900BE3CC051A42198D2834CC690CD0191A6",
            INIT_RAM_1D => X"00936010AD60382DAD58B248C92491101801243002494924A9119A0E8F24B048",
            INIT_RAM_1E => X"4FDA8944931988A494EE44A491FE92491042B5903A016D7EC58824914A491BE9",
            INIT_RAM_1F => X"84A17585424EE150048C92011018036D98F492A414CCC9C1F09CC9AA14926334",
            INIT_RAM_20 => X"4609D8E1DBA440F618F1CC592598D2492CC692193810022A61153761151BBA12",
            INIT_RAM_21 => X"4F3292AB3DEA8DD39D1F853AA6CAF224BD153324B62C7329C2BFF8016D7E1930",
            INIT_RAM_22 => X"BE58EBBE6BBAB81DEEF7F3E72E26522E9650BEC647CF32C64B6C30CF2E4EB9F2",
            INIT_RAM_23 => X"72CF7A7618CE23437AD600F0AC18DE1359762368D31A210E02C2A5D70835DDCC",
            INIT_RAM_24 => X"5AA4D30D6C6B20D4CDAAC045E13C0167BF1A9DA74E8302AAAAAAA1D8A9304A61",
            INIT_RAM_25 => X"48AD62F3C505F4D717EFA505A626B4E9364B3FF75F7DF7DD34193F28B890A630",
            INIT_RAM_26 => X"A93229E53B354935630CB6546EF64A36E677CB6E7D9CCA96A20B56958972B748",
            INIT_RAM_27 => X"FFE007BFEFF247BDF7F03FFC9A48FDE07FF81FF7BFE826C7DBF674F7F2BBB2E8",
            INIT_RAM_28 => X"963BB5DA8001A06D26FB2BA11359AAB6AD5836A0A4E8B0AC2C39140D5D09F83F",
            INIT_RAM_29 => X"2C9242CDBB6D51106D5C6EA8882D1C6EEF64D189573506EDCD982EE62EDD773D",
            INIT_RAM_2A => X"91B09DB6D36F11B198DB8DD8C86DDB6E9B61BB9895035E23E72560CD75FEEBCA",
            INIT_RAM_2B => X"8CF8CB6D69A160B17A04F759864F758C34160A18E272A7F7450C4C47E90C7120",
            INIT_RAM_2C => X"3392B326C2B704AD296AAB2A521E50F2510F25303C87A21710F565F8C77C746F",
            INIT_RAM_2D => X"433AC809B950CEB36AF7F0FA0EB34D8FFEB4AD76EB5632BF7B67ACFF9EF3765D",
            INIT_RAM_2E => X"00000CF191C38D30E60F4EBE8FE6BA1AAA96B5AB6ADBDD6BA5C07A51829B4BF8",
            INIT_RAM_2F => X"3FED978E33FCE79CC1330EC18B653B933B9884609C813F861F771ECCA1B00000",
            INIT_RAM_30 => X"64ACB2FE6D70171D35D5550B43CE7C5B3D93742A17B1887B2CBE7F36E63A5085",
            INIT_RAM_31 => X"2ADF411618B729B83CE1C30096BD63ACC3212F4D17F4B2BE55985573073D11CA",
            INIT_RAM_32 => X"AB48D03D302492491A8DF56BAFD965D19597307EFAA9C7CACB2FA696077F0E83",
            INIT_RAM_33 => X"14D7CB1F4A6D7774DD8810706091577DD4D6B7F4B058594E63FABA74DCB6B3AB",
            INIT_RAM_34 => X"085BCD7B562B99EE579025DD57A0EF64AA69A490F7504C8EB95E5C6768EAD5ED",
            INIT_RAM_35 => X"2A795CD3993DE27B710400000006DE575CD4ABCD3D8BF5A9D9F2DBABDFBC91D9",
            INIT_RAM_36 => X"22A7D89B8BB183BEEEFA3D15DBAE137380BADB29538CA6191867C1C67C1867C7",
            INIT_RAM_37 => X"120006D9BF9A2C9BF619FE17A249AF501CE0148A05C577AF4C794BB386998913",
            INIT_RAM_38 => X"1C15F8798411B2B4575CECC707CCE281B0986F6CE694E717D59BC0B324907F82",
            INIT_RAM_39 => X"2BF9A9F0F9EAB788833D1A6B3DB5706A0F31956BFF97F3A91BBEAED78F45FF22",
            INIT_RAM_3A => X"59588A207921D8C5AB09A6B84AD5B73F000002BD5DE175A687E022B6C0AD4B2B",
            INIT_RAM_3B => X"660CD8C71B3426684B010002013722CA56EF428BA04E7A577B86256FA70374CE",
            INIT_RAM_3C => X"9BD9325D4AEA89F2AEDAD4BBCD350D7F5D769A8B3A6E4761C59005D9D9C9C9E0",
            INIT_RAM_3D => X"BE9BEF4F3EF7EEC93FBB966E9BFAADE507D60EFE6776FFBFF47C1DF78FFEDBFD",
            INIT_RAM_3E => X"EB6BDB7ED9B7AFD7AEAB5AFEA6ECAD66BD72ABD3B8BCEE2F2F6BB59DEEDBF7FB",
            INIT_RAM_3F => X"00005AE23AAE19BA990DCDC5C5E5DAE9935A34D20F6EC8805D59765765DC7B56"
        )
        port map (
            DO => prom_inst_22_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_2,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_23: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0220000000000000080040004023AD496997BBFF877B986EEF16FCF229FA091B",
            INIT_RAM_01 => X"00000000000000000008400000000000000000000000000030600000100007E0",
            INIT_RAM_02 => X"9CDCADCF90E7BD88125BCE706BF6D04AABFC1C001163DC6EFF7FD32303030300",
            INIT_RAM_03 => X"E7622EC485808C841D64B737041FF68813B149A41531A0A612FB14AE2E5B49D4",
            INIT_RAM_04 => X"C52A6A379A382C6D2F5278DA01396D0800C0046405C06F466DD18C4DD7655CD4",
            INIT_RAM_05 => X"AFE59E91BF11498940A0944996D47EE8D7E3A4EAE611AE19A965D01BA86B55E9",
            INIT_RAM_06 => X"042216E0216C85B8912250B7157D5955ADC06CB685BBF071B47D5193363C1CEC",
            INIT_RAM_07 => X"B5D49EA9D7036A45AA9E870B8E8016720C7C3102AE925262492084584942D209",
            INIT_RAM_08 => X"F665955B4E2C63DAC0078652D10120900298F7EE380092442AFD400BEC43C003",
            INIT_RAM_09 => X"D18FCFFFF3FFE7F9FFFFFFF82C0B4221214711E08904524A069491774E663F48",
            INIT_RAM_0A => X"B111114514CB11840E04828849C621392041163C00808D67223422F00110201D",
            INIT_RAM_0B => X"67459F1A8C3240FE4E6A8D028C0C088FCF471D400A11B38211004DD122212288",
            INIT_RAM_0C => X"FE2AC2A884A8CC7FBB821C851CC92B12E15593C0C020FFEE066558590E882D5B",
            INIT_RAM_0D => X"00300A8D128FA20030ACCBAFA237B7024504D36A4BA26081137F059E78991154",
            INIT_RAM_0E => X"09312DACE620656EAF24D57C08FFB14D289613DC32083803B84DC6415FD5EDC0",
            INIT_RAM_0F => X"02E84F961E3C800AC610D276182020227809001A50DDDBA3487BB6AE802BA065",
            INIT_RAM_10 => X"4915C84D6C24BAF53929814CA8A4697E8F4201145AE7415DC122A5F010433107",
            INIT_RAM_11 => X"46AAF6CFDC0791AA97B741995A3B3981E06D1A44D3711955197BB9910FCA2074",
            INIT_RAM_12 => X"3B9254954344968BAC84141C90A9C0E016CB24EDBB4D267E11775FEDD6A2FEB3",
            INIT_RAM_13 => X"0FF81FFF7FFBFFDFFFBFFFE1FF0086F3141AAB6005810C05A1595A893F9D8598",
            INIT_RAM_14 => X"FBFFEFF03FFE0FFFBFAFE0FF80787FFF7FFF83F7F87003FFBFFFFBFFFBFF0FFC",
            INIT_RAM_15 => X"5519198C859000004012AFF4FB060307C92BB732203BFDFEFFFFFFDFFF87FCFF",
            INIT_RAM_16 => X"F40B800FBA159B6DBB296562CB6220EFBE99D2776A202044D9101006FD221D30",
            INIT_RAM_17 => X"1A2955372D510AC266A5445146E27000020C320FAE1557E37154040A10200DC6",
            INIT_RAM_18 => X"111821321BA426A4FE4956B43591D1AC271E83E060341AE5F2023F0808177383",
            INIT_RAM_19 => X"CB9A360865678449975A8AE72B5C0F7BA800C1B5DC55D7D1FE2EF4EED85D00AB",
            INIT_RAM_1A => X"2508062020A0249090009252040249108806A328F4006D2AA514B42FB006ECCC",
            INIT_RAM_1B => X"17C1841358335450D4B26CD2A21B3D8E8211080B81EC040D7FA0B51CD4800811",
            INIT_RAM_1C => X"5B5C1D9D4193E40B9F492B0E0664E13AE35BE6B67AC8057BDACC155F14E906A0",
            INIT_RAM_1D => X"F25E16C87C5D0308EEC52C011514BBC13AFA1028924D0C7CE738105BD47A10AA",
            INIT_RAM_1E => X"1E1EDBBC716D44D2912B80041C44558060CFCC15955C0D600DD5E71393920844",
            INIT_RAM_1F => X"E10F8B8C100323720BEBBDEBB81DF13FF97B252E2CB4F27BA091FBD0002D1A61",
            INIT_RAM_20 => X"DB46809D15D185F8809229B150D05C8081174CA6173B99703DA466629005C604",
            INIT_RAM_21 => X"4EA47F9A7E46083716911B0D585CE937B530218E8D2AD3777EE7D3B4BC56C29A",
            INIT_RAM_22 => X"9434CCA34CC9A1CB1FAACC56168071EAC113F5265D5F6A45A098D604A820508C",
            INIT_RAM_23 => X"538D134115D860ADA57B5B868E54393B1E31E762062577697D57E8464340420E",
            INIT_RAM_24 => X"01859565800698515E10A8189EE9B323E35CE7388D73C6E7A50D0DE6739C73AC",
            INIT_RAM_25 => X"BED23D9A99FF9B77183697955D76BF0CC008822742DA45B88389193DAF094245",
            INIT_RAM_26 => X"00A85E3C5AAE2C49DDC2F6C7B013DACB319A769818A1099A7389F711D76A09BC",
            INIT_RAM_27 => X"A9C9CE3AECF7BE27C000000A8ABA95251B309A60B9DDC19EC3E391458CBB53CA",
            INIT_RAM_28 => X"32EE4CCCECC64F7E6225FC99EC64C3B6DD7DED0FD7CCEA3BF09A006ECDD1009E",
            INIT_RAM_29 => X"D6B97C86DF7D9BEDFB99E36B6658F16C6DEFBDD5DF728D6209C852C37FE67CFF",
            INIT_RAM_2A => X"8662C97BC2E8D3FFDB26D23E87BFD97E635A6560CFD93F8EED26E30C70DE8633",
            INIT_RAM_2B => X"F5569FDE08906765428FB9E6F89FBF0DEAA6064637BCA63FD02E273E5557F054",
            INIT_RAM_2C => X"4EF9AD87727C49CFE7C5DE942B72AC7F6D97DE18920777FDDEE9EB11122A4E18",
            INIT_RAM_2D => X"A1BCE33AD2D8BE40A4E5BB7D7BBEC2CEADBBC8B6F87A4A56FBE0B891DC57E4C6",
            INIT_RAM_2E => X"E0948817C496E9DE8EA1F88F627B7460106691CC4526DCBCCF2CD2F003733C4E",
            INIT_RAM_2F => X"0C840083AD485153ACD3C035591630199B8C096CE4DC557D6D55FCCD738573D6",
            INIT_RAM_30 => X"924C10EFAF3CB9B62486512344C61ADE6F15AB67F335A52513FC85AFAEEE8400",
            INIT_RAM_31 => X"EA4C912568003BB493CE04FF086C188980052BF6ABAAA2FD5D658000011277EB",
            INIT_RAM_32 => X"FFDFFFD75F145247F03A0AE7F1E1EB2D5A99D2444108C6A5CFFD7DEA6ABCC241",
            INIT_RAM_33 => X"02C12B12378356DE2C52041CA7A320C51E0D7CA9F5D575775D57FD75DDFDF75F",
            INIT_RAM_34 => X"6CAFF2622B8D518F63C6030424188FD357718970D25A30CD0731E532DB23002D",
            INIT_RAM_35 => X"D2F8735647315839EF6F683C64773FC73464D5FE354936D50823A5DAEBEBDBCC",
            INIT_RAM_36 => X"59BCEFFBB68A6FF529B3B0D92970010BBB6C7D872421210E190E1CCC47A485EA",
            INIT_RAM_37 => X"5B438D714D4E3DD115E8BD1286EAB5FA1D71BD8F4508BD4BDC8838F9D27B5522",
            INIT_RAM_38 => X"9B96AE83064E84E84C1577BD369FDF5525199894D29B9D3ACCBA3F27D9DC9911",
            INIT_RAM_39 => X"99BA3904854EA910E76808CE76A7998DCB72C49E6429B3F14E73C875B5AE6D35",
            INIT_RAM_3A => X"855EBEA8C1B0000F55D1E716D33CE372B73E6DCF7AD8B2B33111D48F636529AB",
            INIT_RAM_3B => X"800000010000062C649C813BE2639EE988420093314B224ACFFC0FBFFFEA57AB",
            INIT_RAM_3C => X"00000000000000000000000000661EF0F57E0AE0758396AA603052E192CB924D",
            INIT_RAM_3D => X"020028008000524A024A4A284252446240001000101042000054265C7E060000",
            INIT_RAM_3E => X"8004420800620824402040024A1242124204044008404208420A4A42424A1242",
            INIT_RAM_3F => X"990442000864A0284030400454782424440404007E404808A4005448387E547C"
        )
        port map (
            DO => prom_inst_23_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_24: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"B2AA1CB11FBF0000201F8101AF412A8AC5D6525F5C2DD8EF62BAF5B64B7B3199",
            INIT_RAM_01 => X"A41B0424690820860000825904410490DB240E0265A124D018D6D9B8501B9060",
            INIT_RAM_02 => X"8D43C50D9B81601CDE3523D4D0B6984DAD730DA469699B96000B68960874DB50",
            INIT_RAM_03 => X"3AC841F1C073F2A043FDE60C1FEB76A0D07F7C55CBE8112B50A841C1A581A347",
            INIT_RAM_04 => X"476105B47CE4B60006DC8EE263863E89A2E9170FBED2D11EBDB4CEBE2F9D59F6",
            INIT_RAM_05 => X"51CBC8E72C0005404401FFBDDA91816E69BD42CFCAFBABFEB287FE05BE97FCCF",
            INIT_RAM_06 => X"8DB40E7F3C1FC3FAACD555635503F7F8F02DF5D7F6FFCA76EAFDBFF296FABF3E",
            INIT_RAM_07 => X"2032E310821D0A09BFC3F00B171DF5AF7BCE0EF2EA863CF8C002685ABD7CF182",
            INIT_RAM_08 => X"1248A76EFCCAAAA9C6A98E3288AC00828A2003F99FE6DF5A92555FB593A66AC4",
            INIT_RAM_09 => X"A43BD90847E883FFFF7AF2EFD500000015455550555541051415345515F625BB",
            INIT_RAM_0A => X"00287C9742D7BE7F759D999CDC0C0FE896F709DBFFBD3AB7854437749F7D3107",
            INIT_RAM_0B => X"C680989EFC3A06102088AF8F071F7875FF99D11B4A5FFFEE343FDEDDEFE1E7FC",
            INIT_RAM_0C => X"0E755D56FAD6FF7BDCFBF9FF68E6981C8180498C5521DB3311B0D1B3909AD050",
            INIT_RAM_0D => X"0464F37A079D2C9C2E70A38996D1E8A48920C3C33379B288889DA5BE78C6B567",
            INIT_RAM_0E => X"D07B4090C6E9C6DB41A099244653004D4A0B357EF4554441DDDF404451151050",
            INIT_RAM_0F => X"4C0C60613004897FDB9545EDF3716CB6DB561556DB4550E31D55574B72B6DB4C",
            INIT_RAM_10 => X"330FDCCF98101118F475F5F6DB622F7A1CB3FC4E9B019684E020603D998AC161",
            INIT_RAM_11 => X"12B53B6DDB6EDB76DBB6DDB6FFD3F6DF4FB6DDB6EDB76DBF6112678085E4CFC3",
            INIT_RAM_12 => X"70B56CF16772DB6DBB9CE739545FB60459B6587FBDEEDE473330E04043970080",
            INIT_RAM_13 => X"8BA348C33380881206D97AAA2D7CE67776CFF7BDDB8EBF6483C53BAADAAA7E3F",
            INIT_RAM_14 => X"B6DB6DDEE700F73998730C06CEE724EBBC7B0F09DF91C87FE008E60174077610",
            INIT_RAM_15 => X"0410340846EB5D0E04FBB979824A8B700B12B7B1F83C3B067A1B65B6DCDC4E07",
            INIT_RAM_16 => X"431CB2866D1295052166D1399BC9F5BB31315DD71878303A175B8C1C122C71DC",
            INIT_RAM_17 => X"A87CDF5554955100A36C966EF603B75032D972259AD6192893EE9B6581418448",
            INIT_RAM_18 => X"E1334B6105E4296CD683B883900E41B6CB6C31681664F60DEE92AA9331848B7C",
            INIT_RAM_19 => X"DBB6DDB6FB6FFFBDBE6DDBDA965CB7CECDBB0FDAFDFDD5D69BF3F8C75B9D9C5B",
            INIT_RAM_1A => X"B5EEEBDFDCED7B815288F8704C22FF9263CE33B818C620EDB76DBB6DDB6EDB76",
            INIT_RAM_1B => X"796AC79A672F2C253F366B0D9AEAAAEFDFB81FDFFC87F17A19F7F736DB0F012F",
            INIT_RAM_1C => X"99CF45505964498F21E053C2B54A744A3442251BA13B812A82448B0132005A1A",
            INIT_RAM_1D => X"E448E2FAB710EE1862EE72752CD011158A68785808721EDF222A61309B29E84D",
            INIT_RAM_1E => X"0E7038FFB3BF9B8C0AF715197C1AE071FF677EBE5F15EE1E0C3EEEEF7F7777BD",
            INIT_RAM_1F => X"8F9000000FE1B5EA04803821E5518C55AA7211358A5756B89AB0DD53DB4C6C55",
            INIT_RAM_20 => X"B2AA1CB11FBF0000201F8101AF412A8AC5D6525F5C2DD8EF62BAF5B64B7B3199",
            INIT_RAM_21 => X"A41B0424690820860000825904410490DB240E0265A124D018D6D9B8501B9060",
            INIT_RAM_22 => X"8D43C50D9B81601CDE3523D4D0B6984DAD730DA469699B96000B68960874DB50",
            INIT_RAM_23 => X"3AC841F1C073F2A043FDE60C1FEB76A0D07F7C55CBE8112B50A841C1A581A347",
            INIT_RAM_24 => X"476105B47CE4B60006DC8EE263863E89A2E9170FBED2D11EBDB4CEBE2F9D59F6",
            INIT_RAM_25 => X"51CBC8E72C0005404401FFBDDA91816E69BD42CFCAFBABFEB287FE05BE97FCCF",
            INIT_RAM_26 => X"8DB40E7F3C1FC3FAACD555635503F7F8F02DF5D7F6FFCA76EAFDBFF296FABF3E",
            INIT_RAM_27 => X"2032E310821D0A09BFC3F00B171DF5AF7BCE0EF2EA863CF8C002685ABD7CF182",
            INIT_RAM_28 => X"1248A76EFCCAAAA9C6A98E3288AC00828A2003F99FE6DF5A92555FB593A66AC4",
            INIT_RAM_29 => X"A43BD90847E883FFFF7AF2EFD500000015455550555541051415345515F625BB",
            INIT_RAM_2A => X"00287C9742D7BE7F759D999CDC0C0FE896F709DBFFBD3AB7854437749F7D3107",
            INIT_RAM_2B => X"C680989EFC3A06102088AF8F071F7875FF99D11B4A5FFFEE343FDEDDEFE1E7FC",
            INIT_RAM_2C => X"0E755D56FAD6FF7BDCFBF9FF68E6981C8180498C5521DB3311B0D1B3909AD050",
            INIT_RAM_2D => X"0464F37A079D2C9C2E70A38996D1E8A48920C3C33379B288889DA5BE78C6B567",
            INIT_RAM_2E => X"D07B4090C6E9C6DB41A099244653004D4A0B357EF4554441DDDF404451151050",
            INIT_RAM_2F => X"4C0C60613004897FDB9545EDF3716CB6DB561556DB4550E31D55574B72B6DB4C",
            INIT_RAM_30 => X"330FDCCF98101118F475F5F6DB622F7A1CB3FC4E9B019684E020603D998AC161",
            INIT_RAM_31 => X"12B53B6DDB6EDB76DBB6DDB6FFD3F6DF4FB6DDB6EDB76DBF6112678085E4CFC3",
            INIT_RAM_32 => X"70B56CF16772DB6DBB9CE739545FB60459B6587FBDEEDE473330E04043970080",
            INIT_RAM_33 => X"8BA348C33380881206D97AAA2D7CE67776CFF7BDDB8EBF6483C53BAADAAA7E3F",
            INIT_RAM_34 => X"B6DB6DDEE700F73998730C06CEE724EBBC7B0F09DF91C87FE008E60174077610",
            INIT_RAM_35 => X"0410340846EB5D0E04FBB979824A8B700B12B7B1F83C3B067A1B65B6DCDC4E07",
            INIT_RAM_36 => X"431CB2866D1295052166D1399BC9F5BB31315DD71878303A175B8C1C122C71DC",
            INIT_RAM_37 => X"A87CDF5554955100A36C966EF603B75032D972259AD6192893EE9B6581418448",
            INIT_RAM_38 => X"E1334B6105E4296CD683B883900E41B6CB6C31681664F60DEE92AA9331848B7C",
            INIT_RAM_39 => X"DBB6DDB6FB6FFFBDBE6DDBDA965CB7CECDBB0FDAFDFDD5D69BF3F8C75B9D9C5B",
            INIT_RAM_3A => X"B5EEEBDFDCED7B815288F8704C22FF9263CE33B818C620EDB76DBB6DDB6EDB76",
            INIT_RAM_3B => X"796AC79A672F2C253F366B0D9AEAAAEFDFB81FDFFC87F17A19F7F736DB0F012F",
            INIT_RAM_3C => X"99CF45505964498F21E053C2B54A744A3442251BA13B812A82448B0132005A1A",
            INIT_RAM_3D => X"E448E2FAB710EE1862EE72752CD011158A68785808721EDF222A61309B29E84D",
            INIT_RAM_3E => X"0E7038FFB3BF9B8C0AF715197C1AE071FF677EBE5F15EE1E0C3EEEEF7F7777BD",
            INIT_RAM_3F => X"8F9000000FE1B5EA04803821E5518C55AA7211358A5756B89AB0DD53DB4C6C55"
        )
        port map (
            DO => prom_inst_24_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_25: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"B2AA1CB11FBF0000201F8101AF412A8AC5D6525F5C2DD8EF62BAF5B64B7B3199",
            INIT_RAM_01 => X"A41B0424690820860000825904410490DB240E0265A124D018D6D9B8501B9060",
            INIT_RAM_02 => X"8D43C50D9B81601CDE3523D4D0B6984DAD730DA469699B96000B68960874DB50",
            INIT_RAM_03 => X"3AC841F1C073F2A043FDE60C1FEB76A0D07F7C55CBE8112B50A841C1A581A347",
            INIT_RAM_04 => X"476105B47CE4B60006DC8EE263863E89A2E9170FBED2D11EBDB4CEBE2F9D59F6",
            INIT_RAM_05 => X"51CBC8E72C0005404401FFBDDA91816E69BD42CFCAFBABFEB287FE05BE97FCCF",
            INIT_RAM_06 => X"8DB40E7F3C1FC3FAACD555635503F7F8F02DF5D7F6FFCA76EAFDBFF296FABF3E",
            INIT_RAM_07 => X"2032E310821D0A09BFC3F00B171DF5AF7BCE0EF2EA863CF8C002685ABD7CF182",
            INIT_RAM_08 => X"1248A76EFCCAAAA9C6A98E3288AC00828A2003F99FE6DF5A92555FB593A66AC4",
            INIT_RAM_09 => X"A43BD90847E883FFFF7AF2EFD500000015455550555541051415345515F625BB",
            INIT_RAM_0A => X"00287C9742D7BE7F759D999CDC0C0FE896F709DBFFBD3AB7854437749F7D3107",
            INIT_RAM_0B => X"C680989EFC3A06102088AF8F071F7875FF99D11B4A5FFFEE343FDEDDEFE1E7FC",
            INIT_RAM_0C => X"0E755D56FAD6FF7BDCFBF9FF68E6981C8180498C5521DB3311B0D1B3909AD050",
            INIT_RAM_0D => X"0464F37A079D2C9C2E70A38996D1E8A48920C3C33379B288889DA5BE78C6B567",
            INIT_RAM_0E => X"D07B4090C6E9C6DB41A099244653004D4A0B357EF4554441DDDF404451151050",
            INIT_RAM_0F => X"4C0C60613004897FDB9545EDF3716CB6DB561556DB4550E31D55574B72B6DB4C",
            INIT_RAM_10 => X"330FDCCF98101118F475F5F6DB622F7A1CB3FC4E9B019684E020603D998AC161",
            INIT_RAM_11 => X"12B53B6DDB6EDB76DBB6DDB6FFD3F6DF4FB6DDB6EDB76DBF6112678085E4CFC3",
            INIT_RAM_12 => X"70B56CF16772DB6DBB9CE739545FB60459B6587FBDEEDE473330E04043970080",
            INIT_RAM_13 => X"8BA348C33380881206D97AAA2D7CE67776CFF7BDDB8EBF6483C53BAADAAA7E3F",
            INIT_RAM_14 => X"B6DB6DDEE700F73998730C06CEE724EBBC7B0F09DF91C87FE008E60174077610",
            INIT_RAM_15 => X"0410340846EB5D0E04FBB979824A8B700B12B7B1F83C3B067A1B65B6DCDC4E07",
            INIT_RAM_16 => X"431CB2866D1295052166D1399BC9F5BB31315DD71878303A175B8C1C122C71DC",
            INIT_RAM_17 => X"A87CDF5554955100A36C966EF603B75032D972259AD6192893EE9B6581418448",
            INIT_RAM_18 => X"E1334B6105E4296CD683B883900E41B6CB6C31681664F60DEE92AA9331848B7C",
            INIT_RAM_19 => X"DBB6DDB6FB6FFFBDBE6DDBDA965CB7CECDBB0FDAFDFDD5D69BF3F8C75B9D9C5B",
            INIT_RAM_1A => X"B5EEEBDFDCED7B815288F8704C22FF9263CE33B818C620EDB76DBB6DDB6EDB76",
            INIT_RAM_1B => X"796AC79A672F2C253F366B0D9AEAAAEFDFB81FDFFC87F17A19F7F736DB0F012F",
            INIT_RAM_1C => X"99CF45505964498F21E053C2B54A744A3442251BA13B812A82448B0132005A1A",
            INIT_RAM_1D => X"E448E2FAB710EE1862EE72752CD011158A68785808721EDF222A61309B29E84D",
            INIT_RAM_1E => X"0E7038FFB3BF9B8C0AF715197C1AE071FF677EBE5F15EE1E0C3EEEEF7F7777BD",
            INIT_RAM_1F => X"8F9000000FE1B5EA04803821E5518C55AA7211358A5756B89AB0DD53DB4C6C55",
            INIT_RAM_20 => X"B2AA1CB11FBF0000201F8101AF412A8AC5D6525F5C2DD8EF62BAF5B64B7B3199",
            INIT_RAM_21 => X"A41B0424690820860000825904410490DB240E0265A124D018D6D9B8501B9060",
            INIT_RAM_22 => X"8D43C50D9B81601CDE3523D4D0B6984DAD730DA469699B96000B68960874DB50",
            INIT_RAM_23 => X"3AC841F1C073F2A043FDE60C1FEB76A0D07F7C55CBE8112B50A841C1A581A347",
            INIT_RAM_24 => X"476105B47CE4B60006DC8EE263863E89A2E9170FBED2D11EBDB4CEBE2F9D59F6",
            INIT_RAM_25 => X"51CBC8E72C0005404401FFBDDA91816E69BD42CFCAFBABFEB287FE05BE97FCCF",
            INIT_RAM_26 => X"8DB40E7F3C1FC3FAACD555635503F7F8F02DF5D7F6FFCA76EAFDBFF296FABF3E",
            INIT_RAM_27 => X"2032E310821D0A09BFC3F00B171DF5AF7BCE0EF2EA863CF8C002685ABD7CF182",
            INIT_RAM_28 => X"1248A76EFCCAAAA9C6A98E3288AC00828A2003F99FE6DF5A92555FB593A66AC4",
            INIT_RAM_29 => X"A43BD90847E883FFFF7AF2EFD500000015455550555541051415345515F625BB",
            INIT_RAM_2A => X"00287C9742D7BE7F759D999CDC0C0FE896F709DBFFBD3AB7854437749F7D3107",
            INIT_RAM_2B => X"C680989EFC3A06102088AF8F071F7875FF99D11B4A5FFFEE343FDEDDEFE1E7FC",
            INIT_RAM_2C => X"0E755D56FAD6FF7BDCFBF9FF68E6981C8180498C5521DB3311B0D1B3909AD050",
            INIT_RAM_2D => X"0464F37A079D2C9C2E70A38996D1E8A48920C3C33379B288889DA5BE78C6B567",
            INIT_RAM_2E => X"D07B4090C6E9C6DB41A099244653004D4A0B357EF4554441DDDF404451151050",
            INIT_RAM_2F => X"4C0C60613004897FDB9545EDF3716CB6DB561556DB4550E31D55574B72B6DB4C",
            INIT_RAM_30 => X"330FDCCF98101118F475F5F6DB622F7A1CB3FC4E9B019684E020603D998AC161",
            INIT_RAM_31 => X"12B53B6DDB6EDB76DBB6DDB6FFD3F6DF4FB6DDB6EDB76DBF6112678085E4CFC3",
            INIT_RAM_32 => X"70B56CF16772DB6DBB9CE739545FB60459B6587FBDEEDE473330E04043970080",
            INIT_RAM_33 => X"8BA348C33380881206D97AAA2D7CE67776CFF7BDDB8EBF6483C53BAADAAA7E3F",
            INIT_RAM_34 => X"B6DB6DDEE700F73998730C06CEE724EBBC7B0F09DF91C87FE008E60174077610",
            INIT_RAM_35 => X"0410340846EB5D0E04FBB979824A8B700B12B7B1F83C3B067A1B65B6DCDC4E07",
            INIT_RAM_36 => X"431CB2866D1295052166D1399BC9F5BB31315DD71878303A175B8C1C122C71DC",
            INIT_RAM_37 => X"A87CDF5554955100A36C966EF603B75032D972259AD6192893EE9B6581418448",
            INIT_RAM_38 => X"E1334B6105E4296CD683B883900E41B6CB6C31681664F60DEE92AA9331848B7C",
            INIT_RAM_39 => X"DBB6DDB6FB6FFFBDBE6DDBDA965CB7CECDBB0FDAFDFDD5D69BF3F8C75B9D9C5B",
            INIT_RAM_3A => X"B5EEEBDFDCED7B815288F8704C22FF9263CE33B818C620EDB76DBB6DDB6EDB76",
            INIT_RAM_3B => X"796AC79A672F2C253F366B0D9AEAAAEFDFB81FDFFC87F17A19F7F736DB0F012F",
            INIT_RAM_3C => X"99CF45505964498F21E053C2B54A744A3442251BA13B812A82448B0132005A1A",
            INIT_RAM_3D => X"E448E2FAB710EE1862EE72752CD011158A68785808721EDF222A61309B29E84D",
            INIT_RAM_3E => X"0E7038FFB3BF9B8C0AF715197C1AE071FF677EBE5F15EE1E0C3EEEEF7F7777BD",
            INIT_RAM_3F => X"8F9000000FE1B5EA04803821E5518C55AA7211358A5756B89AB0DD53DB4C6C55"
        )
        port map (
            DO => prom_inst_25_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_26: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"1DC952B29949E665F74FDFB109FDBDF6FFAEDDEE62DDDBB1953EC70909090729",
            INIT_RAM_01 => X"80C366581A483526D986E7A412D32E04CC9043233ACDA529DCDF2CB64924B2C9",
            INIT_RAM_02 => X"4612C719B2DDB5ED2F24A636DAD6B660BC19F12641CD62D16326882D8323486D",
            INIT_RAM_03 => X"5FB0371CA3D81111091C3E4081D14471A223DB33046C50B44B3C799660BC81B9",
            INIT_RAM_04 => X"FBFFDDEFF7FFDFDFFEF7FBFDEFFDF54015500EAF933D7F043CF586C8FED5C6FC",
            INIT_RAM_05 => X"9A593E46EBAF66E2DBFAD0001AA56387DDFEFF03F7BDFEDFEDDFDDFFBDFFDEFF",
            INIT_RAM_06 => X"958BBF740E01145450FDC4C3A811F2513E4B24BC7C21659378FBB74F0D10C6FB",
            INIT_RAM_07 => X"78B2D7C3CB9837C620100BC803651CF3F90E34B0FDE20101BC803679CAA3FFFC",
            INIT_RAM_08 => X"0B46E31234F6BB8786BDE4AD66C5AC1B246789C4288D59A110F121304F046688",
            INIT_RAM_09 => X"D35EE96DADB762322222322E9FE780602141399EECE7B5586FAA5F24C6D62066",
            INIT_RAM_0A => X"4E0C19978233336CFFC5B64DDCCC36C376C6FEC5B6DC02EBA5C333870810E231",
            INIT_RAM_0B => X"965303B990C1960F6B2194F66A59A97C749196321E80FB66C45C230DFB2929FC",
            INIT_RAM_0C => X"4E666CA537386E4166C87786CB36479B7CEF32C87F9F32672CA663EC65CE43B5",
            INIT_RAM_0D => X"01400055001007B2C0F87B2F9366C91765334E9DDDF4E32CDB2C53AC894A5B12",
            INIT_RAM_0E => X"180C36FF6E666FCCC32C36CCC1C7FBEBDBB36E75E98060ADB8BA1CA79A300E01",
            INIT_RAM_0F => X"BA9E6F7A581DB36D6E61E6F761BD94BE4DE736DC0B22D86C6464646464666DE1",
            INIT_RAM_10 => X"554015054145104451415541412736DC0B61B61B0D96461774A581C0B6039640",
            INIT_RAM_11 => X"3C78F61C24A81C738843966CC59672AACB2CC000000000000000001555554000",
            INIT_RAM_12 => X"9C0DC40F7DDF0BF786C384C7F09E79E1046E28D8F919F3119BCDE6F3C27E2DDE",
            INIT_RAM_13 => X"0223033980E41856477721B3039EFB37467EF0EE3ECF3DEDBDD6AE7C3ECC2846",
            INIT_RAM_14 => X"C2D926581270ED96C93196191961CBA66E08997099CEC6339D2C88D96032EBB7",
            INIT_RAM_15 => X"F9C0C1C67839F99BA05C607BE8FF1E518679F924BB8B39CE83B75D8C7D6FCDEF",
            INIT_RAM_16 => X"615E40012EE070C3B93E9F90763447004E72641E3463037B38F09A28CF0139EC",
            INIT_RAM_17 => X"C25220467E25A493231980820900008002024012008824080482008491482ED5",
            INIT_RAM_18 => X"F3BF99774CFDD330BAC5A3F6213693B8D7D556DE4FC3333DB63C6C4796D00759",
            INIT_RAM_19 => X"6A565CCF876BE0861ED2DE70000C4266DBCD8B9667BD9D9C99216EB0EE466F72",
            INIT_RAM_1A => X"62692737918D10638E48C6630DB8B1EF6F0FC87BFD3F7AFD89A1C336DFB1230E",
            INIT_RAM_1B => X"EB21253B633F8E0FF79D7258C24448C908806668A035C45C4446DBB318968F4C",
            INIT_RAM_1C => X"6C5E37636CDB6DDA37F3B5AB10E81F01FECF683DB19F5ED8463AF6C7AC929DB1",
            INIT_RAM_1D => X"B6C9B3139866333B9C3CDB6DCDB6DAAAB36DB6E3DB2C6DB6C433B87F5EB06320",
            INIT_RAM_1E => X"77DAEC22DEFECE32C3A33636C28ADB6C9C4E619E3391DCE1E6CE32C3636C28AD",
            INIT_RAM_1F => X"D635F3B9DB7E6E7436DCDB42AAB36F6DBA76DB10D276E6DEF6EEE6988C5BDFDC",
            INIT_RAM_20 => X"F33E75F7A03302261FBB3AFDB6CD9B6DB66CDBBBDA56DB030CE701F4E700E358",
            INIT_RAM_21 => X"F69D8C9284324EC8E498CDC962C8196C840D9B8C933CDB8C46FFF8001FC33B99",
            INIT_RAM_22 => X"D8C3719BB0898BE21FC08D35DCF9B96392C7E46DA6CDDC4304B8685B80D8CB64",
            INIT_RAM_23 => X"D880133F4E790D5AEE66F0660D3EBB7EF08211E046BDE379B98911D14E58479F",
            INIT_RAM_24 => X"281211484D426886D84C8210F49147A505117DA776E16A22222238607CDA635A",
            INIT_RAM_25 => X"368C365C64736B30F396447359C21010000082000400482480251E48C8FE0A85",
            INIT_RAM_26 => X"0F913632D8CB064F0CC27EC3631B39C3B181793B96F366039ECB32037E1D30B6",
            INIT_RAM_27 => X"1FB003FFFBF823FFFFFFC2FE08247EFF8FFFE1FBE000820B27701BCFA6470E38",
            INIT_RAM_28 => X"EBC87239000058364FE890E0E1065F8002C6C3849832C886B5C64B02C6E3F7DF",
            INIT_RAM_29 => X"99659216EDB624F66C8763127B2C8763B5A36C270502C9B7166F638BE377DE77",
            INIT_RAM_2A => X"6EEC36DB6DB5E6E6E76EC37373B765BB6DD86F0332658BCCC1CE997D0F5D573C",
            INIT_RAM_2B => X"23923DB3B679D9CFADEC0CF839C09CDB819D9CF76CAE716192C39771D2C31EDF",
            INIT_RAM_2C => X"115245963609B676E0620B2011812C0DC2C0DCEC226071844C0E189231C91F39",
            INIT_RAM_2D => X"30921610B40C2484D821D09C2484841DEA1B0EB221C887922FC364917867D2C7",
            INIT_RAM_2E => X"0000740CDEB877AEB1A4FDE208CE67E9A48A39A664F3466860238606048C2130",
            INIT_RAM_2F => X"77BD31258739C96196CE43225D1C8E70C7D399187BB4F7664DCED240184C0000",
            INIT_RAM_30 => X"1FC3CE3D9CB0D0FC01CA0443303DE6CA7125B10887A4660669C4CE78CCEFC94C",
            INIT_RAM_31 => X"E0F8B371970E6677F6BC7CDFF228621B1EE1C11879E1381DF877AC50FE440798",
            INIT_RAM_32 => X"8332CC2808D249248778B18300C71CEFBAC50FEA6631307838E3D9C3385A4360",
            INIT_RAM_33 => X"0CDFC01E460412E494560C08112011133CDA2290462626020BAF71DC42030C00",
            INIT_RAM_34 => X"F0F9068DAF94C67330E83045AE1760F6B4E38C30CCFBB3624CC3FC54604831EC",
            INIT_RAM_35 => X"0868206F6EF5BA2700FBFFFFFFF9480709E0009A8C380192C3C0790546676E6E",
            INIT_RAM_36 => X"255C85A7A2C246519956C3BE3322E8DCFA6E5C863E7FFCFFF73EFF33EFF33EFC",
            INIT_RAM_37 => X"02000F890A009F6719E649D18E7AA31231B81E4C8444D19305EFE63DFF628307",
            INIT_RAM_38 => X"E54ABACCF866EDF113F2073C1263496048E415310C0842F9224C441E0000FF02",
            INIT_RAM_39 => X"7EBB5CD134BFBD13C78C08DEC36F389E59870063C951C9FC709A22119A073FD6",
            INIT_RAM_3A => X"78E9C33009CE73C4ECCE9CE6736E721680001170C2E0DCE39CD1666C631BF6DE",
            INIT_RAM_3B => X"2719F7F3C97372E6E7CC555DC888C666646443326731984412498F327900D1CE",
            INIT_RAM_3C => X"E39274C49CE172EA031CC98984D064ED07120804CA4C47894402ACBC47D7D7A0",
            INIT_RAM_3D => X"8E28ED2E7E66D7E49308C1A367680CC26692223C2117EDF339F8047F4CC318EA",
            INIT_RAM_3E => X"25E3EF3F66F38C73E3E318C799658C8E3C12071ACD0EB3434320D2C4626596F0",
            INIT_RAM_3F => X"36DB643FC851E6CE16C8C8C8C8C8F46B4C3811B6CBCF78801C20B2CD2C47CB32"
        )
        port map (
            DO => prom_inst_26_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_2,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_27: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FDDFFFFFFFFFFFFFF7FFBFFFBFDC0A6DBE6F8CFFBB7FEFA39B3DFBF3BEFBB679",
            INIT_RAM_01 => X"FFFFFFFFFFFFFFFFFFF7BFFFFFFFFFFFFFFFFFFFFFFFFFFFCF9FFFFFEFFFF81F",
            INIT_RAM_02 => X"B607E624499300E4DF6D95CB62F62FB75403E400EFBC3BD34080FC9CDCFCFCFF",
            INIT_RAM_03 => X"C9F7627EB100872A52FB5141D65111E6C8DA0ADB6CEC6005C61D0E366B20DCCD",
            INIT_RAM_04 => X"4C3838641E940623ADF28CCA14BCC07104C112BCC9032C48E925594CB886A604",
            INIT_RAM_05 => X"B657485DCD62AC0662C8C005DDE7494C9CA13AAE3234BB0EE1B708A23A2F48AC",
            INIT_RAM_06 => X"96632C3232C3974CDC1172E1779D8C6738251819975DB8146067301E0C0277B6",
            INIT_RAM_07 => X"0776C62C316FF94B0BC3A0288DE6A62B14D6C1A2DADF9BDF85B2CCB02CE1DB2D",
            INIT_RAM_08 => X"07B78D38001FE67E56CCE399DE36D7DDBD699D5CFC5B6D7A1421CE06FE40DB6E",
            INIT_RAM_09 => X"9693E3EFF8FBF1FCEEFBCF7CF9BA6C37640DDF7FFE6187B19ACF089D4C038F66",
            INIT_RAM_0A => X"7CBBCB2CB384BD0D92ED105D0617856E80441124B31DE58B8C001607FEE66889",
            INIT_RAM_0B => X"3D3CF1BE8C84DDB000565880A776E5C0E13166E49F47119A4CA1311CF97B965E",
            INIT_RAM_0C => X"7EE296E8986E64C6DCDDE59436641567648CB84DEB7D7937F974F038D838274F",
            INIT_RAM_0D => X"1889D25CB816ACC6627802052C61A4099B7B0EC923971DB3B9F9204BDBCCFA45",
            INIT_RAM_0E => X"7D361CDE72B925658DBE1F7C4707E195C5C665B8118C3C31B196C261DA85A5E1",
            INIT_RAM_0F => X"1C5CF062CA6F13854A59BDEEEA07E3C6559EBB3618111895CBBACCBCD512B5F0",
            INIT_RAM_10 => X"2EB0B348C0B62337739B1BC73192392592C84E37B7AC141CFE65EE76D83CB083",
            INIT_RAM_11 => X"1D77401A0C0CCF5DEEE561F7F7E68CBE72E48E570B047C772CBACC33753080E3",
            INIT_RAM_12 => X"19B9466E6D7B527565924244B20C5DA22B60D21B6030D9960699E11209699604",
            INIT_RAM_13 => X"F7F7FDDFFEDFF6FF7FFEEFFEFEFC4E51EC0888848E1F2246347B66608D8A3B39",
            INIT_RAM_14 => X"FFDFFF6FFFBDFFDFFF57FF7F7FB7FBBDFBDFFDBFF78FFDBFFEDDFFFDFFFEFF6F",
            INIT_RAM_15 => X"CEEC06DAECB0001569589D5F267AFE086C8FED5DE41DFEFF027DFDFF7FFBFBFD",
            INIT_RAM_16 => X"BA42813453FF4EDB60C6BF8DB6E267BC56CB69BBCE636CCCB3B2B4B103CC46D5",
            INIT_RAM_17 => X"881331ED7AC4EFD38DFACDBB236790005719AEA2FAECCF0D126A30A27562C61B",
            INIT_RAM_18 => X"CE618EEDCFB393738178C476C36CB61F71307F6803F677575763DB2D8C3118E4",
            INIT_RAM_19 => X"36DB5B7BD2850018CF936621C6863095A73F7BE7442CB13310B9C0BBB96EEF16",
            INIT_RAM_1A => X"0408002024010408824080002008091482ED5615E40012EE630C3B2CDB2C13A7",
            INIT_RAM_1B => X"4A3E508B49DC6BEAAB4F3F0CCCF6D8F468F2DA00EB384A7F5324932319800010",
            INIT_RAM_1C => X"2E43664448EFF19872648DBACEEDB76E26439BCCEF2DFBF664594B04FBAE72A8",
            INIT_RAM_1D => X"3DA139003D7A86B2F878DD99DAFB70DE1A19F3FB7DB3B8EF2633007664CB1999",
            INIT_RAM_1E => X"EFF4FDE394D0E19B6FD89186C23CF071E6F1CC8F7FC4F1E48756B0DCD8ED6D0C",
            INIT_RAM_1F => X"3C766E63DB6481CB39BC8C68831C724633186CC1BAE9D608A5DEF0FF219C28C1",
            INIT_RAM_20 => X"24C921BB3332DC66D9C1706B6C5903129639A3BA4088EDB496EDBBBFC2CC40B6",
            INIT_RAM_21 => X"FF7CCCEFE1996DE3ED6D8CFBF1871BD98EE7646242664EB2E338BD0098386371",
            INIT_RAM_22 => X"63FC93ED92CA4DC61B01639318985C88F01680E307C42311C0124700B28BF9B4",
            INIT_RAM_23 => X"414D536A41D144B6C4624A2B00366D8CF6734A4A2DC465B308462CCBD1BF9CB8",
            INIT_RAM_24 => X"CB76E03779E019E2C4E4028219C38C202C9384E0D24E569C2E4D4D60B670CE37",
            INIT_RAM_25 => X"E1265727652C8F0C422BA8C28A0FBB893B0881E00403DDD8843B2D8EB929D0D8",
            INIT_RAM_26 => X"C228A2050470925E29A35D8D06242712CD25C924189820CD85A710947C802013",
            INIT_RAM_27 => X"5F9CB25A3631964C20007FF5754FC631A97D4F93986C30CF24394625658DE9A7",
            INIT_RAM_28 => X"C7E1B221EA10E38F64EF31CEBF3368E1C712BB1B33781134CFE54C2123349A6E",
            INIT_RAM_29 => X"7DCCFC5939C4EC79CF0E1CD43BA7AFC716900A21BDB9DD0FCC7ECE1063238407",
            INIT_RAM_2A => X"499D7BD86619EE5574CD27C80D39F71E653FDCF1B366737233CBB98D1E7B330F",
            INIT_RAM_2B => X"AAAD6B6AF36195DA637C6EFA3E36E8FE97FA02EC26EB46198AD8DAD8C11260AF",
            INIT_RAM_2C => X"C23B9D130CA49818913D3A2C1FBF71C5B0C774336F903C677D976189D98CA127",
            INIT_RAM_2D => X"CEC3000F432029B3FE3F211712944CA54D1940F193204C199C9F49666BC11B38",
            INIT_RAM_2E => X"2F3982C7BE09AD4A32196807648A2495ADF98FD2B15E604B52F12FBBC811C953",
            INIT_RAM_2F => X"E33CB578DEBFAFAEDFD530DE8FA1992072F31B116644B18C72F9F44116C79ADF",
            INIT_RAM_30 => X"7FB1E62675F7C2CBE01032DCA16BADC570C1CBF7ECBC4E7E6C5425D4550BE1A8",
            INIT_RAM_31 => X"59F878FCF5689FCFEF34BFD52FA2422A56A3C113409F7813007F8D6B5F80FE9D",
            INIT_RAM_32 => X"00000008800AC11D556264251ECFA68C056FBCCB040C614A0240000300D2F6FF",
            INIT_RAM_33 => X"C744FD00E1A7F9E9FBFE4777FD50ABD11F0E57FF4808802282200888A20AA880",
            INIT_RAM_34 => X"57781E91788044213E091339886F337D0612CA646CD48FC58EE77EDD7ECEC466",
            INIT_RAM_35 => X"662FF5DF9CB107BB23A39EF7B95E7372200448DBDC18F9C0DE0EF379BF494806",
            INIT_RAM_36 => X"06F6612D770080980A40D293FEC069F16CB2164CA033C539F69B37741AEF1CE3",
            INIT_RAM_37 => X"0100046606572583002086010800054C0F2DE8371AC0000A9003E024840C7C08",
            INIT_RAM_38 => X"8461D33183C33C33D27577FCFE7FCF2572CBE0000C02060C000C0DF50F68A580",
            INIT_RAM_39 => X"9EC30492764D54DF999727A18953C642308C32411294092663883EC848622649",
            INIT_RAM_3A => X"81102007A7C0000B18CF6AC83C9B581F9891332601CE48E34EFBC607389C5D55",
            INIT_RAM_3B => X"800000007FFCEC621355B688B1D849BB6608185970D976205800000000070103",
            INIT_RAM_3C => X"00000000000000000000000000005290977202A255393471055CA904CBAE2493",
            INIT_RAM_3D => X"0400000000000C34023C2E302464003C00000000000000000020460024000000",
            INIT_RAM_3E => X"80084204004204423E1E3E02247E3C7E3C7E7E7E7E30007E3C7E7E7E3C7E7C3C",
            INIT_RAM_3F => X"4200420000441C443C0C3C00480018FC387C7C000000007E1800383000002048"
        )
        port map (
            DO => prom_inst_27_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_28: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"34AE14114000000000000001AC042A88C586125F1C3418006280F5804B790391",
            INIT_RAM_01 => X"80194E74210820060001864B4D0082080021270865A1259019925CB0C01BA070",
            INIT_RAM_02 => X"9F43CD0D8F01601CDE1523F450B2884CAD6304AC2B68BBB28A1B29B29865D950",
            INIT_RAM_03 => X"1EC8C1F9C07AF00243F5A5F40BEB5A90E03F3E0CC3A42121000840C08581A107",
            INIT_RAM_04 => X"676385B45DE23A8006D68480C1043A9AA1E0171E187AD1169EF458BE2F9C1196",
            INIT_RAM_05 => X"30CB4AFF2C00554401140129511181606BBC48CFCAF2ABD83087FE249497F647",
            INIT_RAM_06 => X"8EF400000000000804D999BD00000000B124A417FE5FD2526AFF97F4925ABF36",
            INIT_RAM_07 => X"303A6311821D0C0936A1C00A023DCF077ADE1AF3E8865CE8C082785C1F6CD183",
            INIT_RAM_08 => X"1089067CA8EAAAA806A8163308A601861A6003F91FE75BDADB55500E8286AAC4",
            INIT_RAM_09 => X"802B5C1C468062FDD77A7ABFC5000000155555541555050514402455150F2692",
            INIT_RAM_0A => X"40282A56A2D5BED2D59A444D9BDA1F803A730BC9ABAD2AB3880415548B357003",
            INIT_RAM_0B => X"CF8089C8989A04301E982FA902335435FB8B00C95A4FFAA7302ADA48EFA1FDAC",
            INIT_RAM_0C => X"0E344E46BAC2B000020009DA60EE8809A10849AE5145D9B60090D11B15DA10D0",
            INIT_RAM_0D => X"5524B1DE058D2C9C2EF0A38196C5E8AD8B024100318B368888B001BEF8C6B422",
            INIT_RAM_0E => X"F07900848240824942009130525700474C09603E74174441C88B405141541410",
            INIT_RAM_0F => X"0424352170000132499544A4D9392D9249523552494FF0E10555540932924C08",
            INIT_RAM_10 => X"1107DDDF98303139FC7CFCF2493C26905D90044A13011208E060603D99F2CE61",
            INIT_RAM_11 => X"16B59924C926493249924C9271D7F24F4F924C926493249F63B2EF81C5E447E3",
            INIT_RAM_12 => X"6009EC1126765924994A5299544C92084BB2487DF56E4E47311060C0C1B34180",
            INIT_RAM_13 => X"8AE1C9431180891004D982AA257CE23712DFBEADC98EBF6483DD2B4BDAAA073D",
            INIT_RAM_14 => X"B2C924DCE7008432887304166E6365F99C5A0B19CE98D83BE088E0017C077633",
            INIT_RAM_15 => X"0410240904AA190608921BFB864C995143131DE39ABC1B023A0B24925E4C4692",
            INIT_RAM_16 => X"410C9282651290002164F17D9BEDF0211E714C920938305B0553CC0C32443354",
            INIT_RAM_17 => X"E83CD004029C1700E03DB366F20A9392764D722D8E561928B36E992581418448",
            INIT_RAM_18 => X"033BF36301E2012ED281B883B406C096492C11293664F604E790AAB3318C8B20",
            INIT_RAM_19 => X"49924C927B2F94D49B25CBDF861A93CE49932BCAFFC7F5E919C128C249DEBC1B",
            INIT_RAM_1A => X"D5A4CEFB4CF569C15384F4F0CA62FF9653D936F8094A40E493249924C9264932",
            INIT_RAM_1B => X"FAEBEFB6F7555D6DBD762B1D8AFFEA00000000000C83712E01BED332490D820F",
            INIT_RAM_1C => X"B95E445DFAED5BABF5E56BCAF49A7CD228D2A8DB895B896288C990CBB212D21A",
            INIT_RAM_1D => X"C44C80FAB7006E19E26E00652DC21140032858F808720A55202AC160BB29684C",
            INIT_RAM_1E => X"0E3030BA929B8BA40A773F192812E06175253EBE5F15E61A249E6667382223BC",
            INIT_RAM_1F => X"8F9000000FB5D5E600901221E9700C55AA0631E10B5E04A890204D504946ECFD",
            INIT_RAM_20 => X"34AE14114000000000000001AC042A88C586125F1C3418006280F5804B790391",
            INIT_RAM_21 => X"80194E74210820060001864B4D0082080021270865A1259019925CB0C01BA070",
            INIT_RAM_22 => X"9F43CD0D8F01601CDE1523F450B2884CAD6304AC2B68BBB28A1B29B29865D950",
            INIT_RAM_23 => X"1EC8C1F9C07AF00243F5A5F40BEB5A90E03F3E0CC3A42121000840C08581A107",
            INIT_RAM_24 => X"676385B45DE23A8006D68480C1043A9AA1E0171E187AD1169EF458BE2F9C1196",
            INIT_RAM_25 => X"30CB4AFF2C00554401140129511181606BBC48CFCAF2ABD83087FE249497F647",
            INIT_RAM_26 => X"8EF400000000000804D999BD00000000B124A417FE5FD2526AFF97F4925ABF36",
            INIT_RAM_27 => X"303A6311821D0C0936A1C00A023DCF077ADE1AF3E8865CE8C082785C1F6CD183",
            INIT_RAM_28 => X"1089067CA8EAAAA806A8163308A601861A6003F91FE75BDADB55500E8286AAC4",
            INIT_RAM_29 => X"802B5C1C468062FDD77A7ABFC5000000155555541555050514402455150F2692",
            INIT_RAM_2A => X"40282A56A2D5BED2D59A444D9BDA1F803A730BC9ABAD2AB3880415548B357003",
            INIT_RAM_2B => X"CF8089C8989A04301E982FA902335435FB8B00C95A4FFAA7302ADA48EFA1FDAC",
            INIT_RAM_2C => X"0E344E46BAC2B000020009DA60EE8809A10849AE5145D9B60090D11B15DA10D0",
            INIT_RAM_2D => X"5524B1DE058D2C9C2EF0A38196C5E8AD8B024100318B368888B001BEF8C6B422",
            INIT_RAM_2E => X"F07900848240824942009130525700474C09603E74174441C88B405141541410",
            INIT_RAM_2F => X"0424352170000132499544A4D9392D9249523552494FF0E10555540932924C08",
            INIT_RAM_30 => X"1107DDDF98303139FC7CFCF2493C26905D90044A13011208E060603D99F2CE61",
            INIT_RAM_31 => X"16B59924C926493249924C9271D7F24F4F924C926493249F63B2EF81C5E447E3",
            INIT_RAM_32 => X"6009EC1126765924994A5299544C92084BB2487DF56E4E47311060C0C1B34180",
            INIT_RAM_33 => X"8AE1C9431180891004D982AA257CE23712DFBEADC98EBF6483DD2B4BDAAA073D",
            INIT_RAM_34 => X"B2C924DCE7008432887304166E6365F99C5A0B19CE98D83BE088E0017C077633",
            INIT_RAM_35 => X"0410240904AA190608921BFB864C995143131DE39ABC1B023A0B24925E4C4692",
            INIT_RAM_36 => X"410C9282651290002164F17D9BEDF0211E714C920938305B0553CC0C32443354",
            INIT_RAM_37 => X"E83CD004029C1700E03DB366F20A9392764D722D8E561928B36E992581418448",
            INIT_RAM_38 => X"033BF36301E2012ED281B883B406C096492C11293664F604E790AAB3318C8B20",
            INIT_RAM_39 => X"49924C927B2F94D49B25CBDF861A93CE49932BCAFFC7F5E919C128C249DEBC1B",
            INIT_RAM_3A => X"D5A4CEFB4CF569C15384F4F0CA62FF9653D936F8094A40E493249924C9264932",
            INIT_RAM_3B => X"FAEBEFB6F7555D6DBD762B1D8AFFEA00000000000C83712E01BED332490D820F",
            INIT_RAM_3C => X"B95E445DFAED5BABF5E56BCAF49A7CD228D2A8DB895B896288C990CBB212D21A",
            INIT_RAM_3D => X"C44C80FAB7006E19E26E00652DC21140032858F808720A55202AC160BB29684C",
            INIT_RAM_3E => X"0E3030BA929B8BA40A773F192812E06175253EBE5F15E61A249E6667382223BC",
            INIT_RAM_3F => X"8F9000000FB5D5E600901221E9700C55AA0631E10B5E04A890204D504946ECFD"
        )
        port map (
            DO => prom_inst_28_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_29: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"34AE14114000000000000001AC042A88C586125F1C3418006280F5804B790391",
            INIT_RAM_01 => X"80194E74210820060001864B4D0082080021270865A1259019925CB0C01BA070",
            INIT_RAM_02 => X"9F43CD0D8F01601CDE1523F450B2884CAD6304AC2B68BBB28A1B29B29865D950",
            INIT_RAM_03 => X"1EC8C1F9C07AF00243F5A5F40BEB5A90E03F3E0CC3A42121000840C08581A107",
            INIT_RAM_04 => X"676385B45DE23A8006D68480C1043A9AA1E0171E187AD1169EF458BE2F9C1196",
            INIT_RAM_05 => X"30CB4AFF2C00554401140129511181606BBC48CFCAF2ABD83087FE249497F647",
            INIT_RAM_06 => X"8EF400000000000804D999BD00000000B124A417FE5FD2526AFF97F4925ABF36",
            INIT_RAM_07 => X"303A6311821D0C0936A1C00A023DCF077ADE1AF3E8865CE8C082785C1F6CD183",
            INIT_RAM_08 => X"1089067CA8EAAAA806A8163308A601861A6003F91FE75BDADB55500E8286AAC4",
            INIT_RAM_09 => X"802B5C1C468062FDD77A7ABFC5000000155555541555050514402455150F2692",
            INIT_RAM_0A => X"40282A56A2D5BED2D59A444D9BDA1F803A730BC9ABAD2AB3880415548B357003",
            INIT_RAM_0B => X"CF8089C8989A04301E982FA902335435FB8B00C95A4FFAA7302ADA48EFA1FDAC",
            INIT_RAM_0C => X"0E344E46BAC2B000020009DA60EE8809A10849AE5145D9B60090D11B15DA10D0",
            INIT_RAM_0D => X"5524B1DE058D2C9C2EF0A38196C5E8AD8B024100318B368888B001BEF8C6B422",
            INIT_RAM_0E => X"F07900848240824942009130525700474C09603E74174441C88B405141541410",
            INIT_RAM_0F => X"0424352170000132499544A4D9392D9249523552494FF0E10555540932924C08",
            INIT_RAM_10 => X"1107DDDF98303139FC7CFCF2493C26905D90044A13011208E060603D99F2CE61",
            INIT_RAM_11 => X"16B59924C926493249924C9271D7F24F4F924C926493249F63B2EF81C5E447E3",
            INIT_RAM_12 => X"6009EC1126765924994A5299544C92084BB2487DF56E4E47311060C0C1B34180",
            INIT_RAM_13 => X"8AE1C9431180891004D982AA257CE23712DFBEADC98EBF6483DD2B4BDAAA073D",
            INIT_RAM_14 => X"B2C924DCE7008432887304166E6365F99C5A0B19CE98D83BE088E0017C077633",
            INIT_RAM_15 => X"0410240904AA190608921BFB864C995143131DE39ABC1B023A0B24925E4C4692",
            INIT_RAM_16 => X"410C9282651290002164F17D9BEDF0211E714C920938305B0553CC0C32443354",
            INIT_RAM_17 => X"E83CD004029C1700E03DB366F20A9392764D722D8E561928B36E992581418448",
            INIT_RAM_18 => X"033BF36301E2012ED281B883B406C096492C11293664F604E790AAB3318C8B20",
            INIT_RAM_19 => X"49924C927B2F94D49B25CBDF861A93CE49932BCAFFC7F5E919C128C249DEBC1B",
            INIT_RAM_1A => X"D5A4CEFB4CF569C15384F4F0CA62FF9653D936F8094A40E493249924C9264932",
            INIT_RAM_1B => X"FAEBEFB6F7555D6DBD762B1D8AFFEA00000000000C83712E01BED332490D820F",
            INIT_RAM_1C => X"B95E445DFAED5BABF5E56BCAF49A7CD228D2A8DB895B896288C990CBB212D21A",
            INIT_RAM_1D => X"C44C80FAB7006E19E26E00652DC21140032858F808720A55202AC160BB29684C",
            INIT_RAM_1E => X"0E3030BA929B8BA40A773F192812E06175253EBE5F15E61A249E6667382223BC",
            INIT_RAM_1F => X"8F9000000FB5D5E600901221E9700C55AA0631E10B5E04A890204D504946ECFD",
            INIT_RAM_20 => X"34AE14114000000000000001AC042A88C586125F1C3418006280F5804B790391",
            INIT_RAM_21 => X"80194E74210820060001864B4D0082080021270865A1259019925CB0C01BA070",
            INIT_RAM_22 => X"9F43CD0D8F01601CDE1523F450B2884CAD6304AC2B68BBB28A1B29B29865D950",
            INIT_RAM_23 => X"1EC8C1F9C07AF00243F5A5F40BEB5A90E03F3E0CC3A42121000840C08581A107",
            INIT_RAM_24 => X"676385B45DE23A8006D68480C1043A9AA1E0171E187AD1169EF458BE2F9C1196",
            INIT_RAM_25 => X"30CB4AFF2C00554401140129511181606BBC48CFCAF2ABD83087FE249497F647",
            INIT_RAM_26 => X"8EF400000000000804D999BD00000000B124A417FE5FD2526AFF97F4925ABF36",
            INIT_RAM_27 => X"303A6311821D0C0936A1C00A023DCF077ADE1AF3E8865CE8C082785C1F6CD183",
            INIT_RAM_28 => X"1089067CA8EAAAA806A8163308A601861A6003F91FE75BDADB55500E8286AAC4",
            INIT_RAM_29 => X"802B5C1C468062FDD77A7ABFC5000000155555541555050514402455150F2692",
            INIT_RAM_2A => X"40282A56A2D5BED2D59A444D9BDA1F803A730BC9ABAD2AB3880415548B357003",
            INIT_RAM_2B => X"CF8089C8989A04301E982FA902335435FB8B00C95A4FFAA7302ADA48EFA1FDAC",
            INIT_RAM_2C => X"0E344E46BAC2B000020009DA60EE8809A10849AE5145D9B60090D11B15DA10D0",
            INIT_RAM_2D => X"5524B1DE058D2C9C2EF0A38196C5E8AD8B024100318B368888B001BEF8C6B422",
            INIT_RAM_2E => X"F07900848240824942009130525700474C09603E74174441C88B405141541410",
            INIT_RAM_2F => X"0424352170000132499544A4D9392D9249523552494FF0E10555540932924C08",
            INIT_RAM_30 => X"1107DDDF98303139FC7CFCF2493C26905D90044A13011208E060603D99F2CE61",
            INIT_RAM_31 => X"16B59924C926493249924C9271D7F24F4F924C926493249F63B2EF81C5E447E3",
            INIT_RAM_32 => X"6009EC1126765924994A5299544C92084BB2487DF56E4E47311060C0C1B34180",
            INIT_RAM_33 => X"8AE1C9431180891004D982AA257CE23712DFBEADC98EBF6483DD2B4BDAAA073D",
            INIT_RAM_34 => X"B2C924DCE7008432887304166E6365F99C5A0B19CE98D83BE088E0017C077633",
            INIT_RAM_35 => X"0410240904AA190608921BFB864C995143131DE39ABC1B023A0B24925E4C4692",
            INIT_RAM_36 => X"410C9282651290002164F17D9BEDF0211E714C920938305B0553CC0C32443354",
            INIT_RAM_37 => X"E83CD004029C1700E03DB366F20A9392764D722D8E561928B36E992581418448",
            INIT_RAM_38 => X"033BF36301E2012ED281B883B406C096492C11293664F604E790AAB3318C8B20",
            INIT_RAM_39 => X"49924C927B2F94D49B25CBDF861A93CE49932BCAFFC7F5E919C128C249DEBC1B",
            INIT_RAM_3A => X"D5A4CEFB4CF569C15384F4F0CA62FF9653D936F8094A40E493249924C9264932",
            INIT_RAM_3B => X"FAEBEFB6F7555D6DBD762B1D8AFFEA00000000000C83712E01BED332490D820F",
            INIT_RAM_3C => X"B95E445DFAED5BABF5E56BCAF49A7CD228D2A8DB895B896288C990CBB212D21A",
            INIT_RAM_3D => X"C44C80FAB7006E19E26E00652DC21140032858F808720A55202AC160BB29684C",
            INIT_RAM_3E => X"0E3030BA929B8BA40A773F192812E06175253EBE5F15E61A249E6667382223BC",
            INIT_RAM_3F => X"8F9000000FB5D5E600901221E9700C55AA0631E10B5E04A890204D504946ECFD"
        )
        port map (
            DO => prom_inst_29_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_30: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0C454AE52948A455454D1E1109D431C4FA28598C0250EB311118030909090741",
            INIT_RAM_01 => X"10080078412401200206C59008402692C4484322BA442C00C45B2DB6C96592CB",
            INIT_RAM_02 => X"CC16830D90DDB9810F6DA616DAD6B6D21819C32E40A56241233780AD03242400",
            INIT_RAM_03 => X"88903C5CE1001110190C2244A0800451A222D9B6002440942911648A501881B4",
            INIT_RAM_04 => X"0004000080080001000080200040000015555C0630313104304492D84A150644",
            INIT_RAM_05 => X"8881B84EEB2C022201A3500020294BA750000001000020020001000400020001",
            INIT_RAM_06 => X"55AA0770101101444488C4628232165122C364A05C6461B3789A345C0D30C471",
            INIT_RAM_07 => X"38E213078980478061301ED00B3505B6FA1A351829621100ED00B6DB4EA68BD4",
            INIT_RAM_08 => X"8900E71414778B86C095A2AD6706902024420100288D59A1201163045C048088",
            INIT_RAM_09 => X"D38EE864A49362322222322E9FE4806001C479BC6DE7B57067C243270612A182",
            INIT_RAM_0A => X"460C18B3C2333360004D96CCCDC4324332427C44925C02EB214611831810E238",
            INIT_RAM_0B => X"9251233C92449706212094734A51AB7CE091B6761E80F926C04C2204FE21297A",
            INIT_RAM_0C => X"CE6C64A432106441464432424A3205193DCE00887F9F332728C643EC64844110",
            INIT_RAM_0D => X"01D000555515571240F8796796265B1725160E9CC0C4E22C59240104894C59B6",
            INIT_RAM_0E => X"1018627F2664278C4364324440C6BBB9D9126424C10842A490A848F29A001C01",
            INIT_RAM_0F => X"901B2630481C93272621E3E2219DA53B04E3324A0926C864ECECECECECEE25F1",
            INIT_RAM_10 => X"5540005540150541451044510163324A092192190CB24C32600481C19203B220",
            INIT_RAM_11 => X"3060C60C24280C330041B2658CBF36AE597E4000000000000000000000001555",
            INIT_RAM_12 => X"900504140DCF8A3208040C484188688304803801A301C1120904824106F86F18",
            INIT_RAM_13 => X"0464033980E42006CFC7003105BEF373A008C0803001102C07120A30220C0088",
            INIT_RAM_14 => X"024B6E60966084B25B71981B1980CA0C2408B9419BCE4211080C9818607283F7",
            INIT_RAM_15 => X"E0E0E2023A993189A04CA03BF8FF08808639E8649B9B38EE843F4C90512504A1",
            INIT_RAM_16 => X"0020BFFFFEA08043A9001FB0769C4B005A726C1E9C65037968509A484F413B3C",
            INIT_RAM_17 => X"004268D66A24A497005D80820100480022000902408000802090448080400000",
            INIT_RAM_18 => X"733301605EF817B14005B3E6633290208085F09EC61010040610CCC79EC08540",
            INIT_RAM_19 => X"6AD61DCC0409018E1010DE400000C666CB0C0396661011BBC4937892CECEE736",
            INIT_RAM_1A => X"06696577118D10238E58C7631DB833E4470BC831C51E397A98D0C01603526106",
            INIT_RAM_1B => X"A52325352162180DF0B4B2D8C244484908807778A00104104444498101938104",
            INIT_RAM_1C => X"222D3721264924DE07C3B1AB30EA1C01EA1C40BA90912D4840296A4295B29A91",
            INIT_RAM_1D => X"9245EB108C06332E0C1CE925C4924AAAD924938B992424924C33B8EFAE90EA94",
            INIT_RAM_1E => X"435AE46248F8C61243E4B212471649245C42301E33917060E746124B21243164",
            INIT_RAM_1F => X"5214B28089362024125C4942AAD92724B9764930D24550D8568D50988C491F1C",
            INIT_RAM_20 => X"C3785AF7A012816618F5AD7C92C6C924963649BB92424B012C02007402002148",
            INIT_RAM_21 => X"C6B99CB78476DE58E5B8DDDB62481B64840C954493381544C0FFF80113633B9B",
            INIT_RAM_22 => X"D8C3588AF9999BE0175227341DE039E193C3E82626CD10410CEC041B41D8C36E",
            INIT_RAM_23 => X"4988133D0C681F0246661E2D0C3899FB108191A1409CE30D949B31515E5C47D6",
            INIT_RAM_24 => X"3820130044026704C0088008D2510FE7071075A542F12000000009200CCE2658",
            INIT_RAM_25 => X"168C1E4824294971F38604294B0258300006096412DB6C94924800682F351CA4",
            INIT_RAM_26 => X"0FB434326C5F06CF1CC625C363BB1913B180591B1251660182593201882030B2",
            INIT_RAM_27 => X"0000062008000621040402000000C00808020100200010096F521BCF8E4F0E38",
            INIT_RAM_28 => X"FB78F2790000C8324EE890C08102FF8247C381848036C8879582C907C6470000",
            INIT_RAM_29 => X"99249016CDB62C12E487631609648763B5A3246304024BB6162FE30BE367CAF7",
            INIT_RAM_2A => X"6EEC365B65B9A6C4E66EC362733665B32DD86D022A61D34E418A98781E0D031D",
            INIT_RAM_2B => X"21921C9792F8994F8DFC1CF878818CD3108994E624CE7260B2479B32D6470EDF",
            INIT_RAM_2C => X"00D245961E019272600007203083241CC241CCEC2220F184441E489210C90E19",
            INIT_RAM_2D => X"1092161134042485F842D0AC2485A49BA0134C1220CD87942563E4A128677242",
            INIT_RAM_2E => X"000070184C98F3A6B1E5F38608CEEFB9048C290644B24A40E0230E0C04052170",
            INIT_RAM_2F => X"F69D31248F39C923B2D9C362CD8E9620C5939B183BBCF7260A5ED640085C0000",
            INIT_RAM_30 => X"1CC1C65DBCB0C1FC10CF0442107DE7CA712DB10885A4220EE9C4CE78CDEFC98C",
            INIT_RAM_31 => X"A0B093709616E6F7F2BC7CFDF220423936E1E34C1BE1281CF8330C40FE4D01B8",
            INIT_RAM_32 => X"0232CC00080000048F7CF18280E38CE7D0C40FC06231304C1C65DBC33A59C361",
            INIT_RAM_33 => X"245D420AC0063B74B092240811221111145EB0D846262E020A6F59DC42130D01",
            INIT_RAM_34 => X"C0FD86A6AD80C2B33AE81084A63370F395E79E70EEF903640CEBD434C05870A9",
            INIT_RAM_35 => X"0048302E6EE1380E2104210888096C0789E8419F9E18011766E02D030B676EAE",
            INIT_RAM_36 => X"015885A5A6424651995383BE732381C8FE0610003EC7FD8FF62EFF62EFF22EFC",
            INIT_RAM_37 => X"02000F8012081F7681E619D38EFAA71231983E2584C4138345E6A63D9F720205",
            INIT_RAM_38 => X"6940195AE006B03116110C360AD38920486415009D0000F12028C21E0001FE02",
            INIT_RAM_39 => X"08180AF134F8B119C3842818003118182B4400C11B518B8C410A22111E043FCA",
            INIT_RAM_3A => X"F8F9C1703B5C9448C5A63C4D316AE00480001131C2A08C719C916630E00C4018",
            INIT_RAM_3B => X"2008F3E82932AA6557C055539C49C616E4624764E333184C22419B22EC01F1DE",
            INIT_RAM_3C => X"729A51E694B1734B0310E3CD06182CC9879B0C05886045008202AC9C82C282E0",
            INIT_RAM_3D => X"1431493AEB4C93649308C1A22E4C0E8274B024582224C93559D008A668939142",
            INIT_RAM_3E => X"35B3ADBD66DB08FB73721084C9768E9B3E13031A4D0E93434330DA4467650C21",
            INIT_RAM_3F => X"00006E3FC804E6CE0248C8C8C8C8F54B4828503A4F0738801820BB47B488439B"
        )
        port map (
            DO => prom_inst_30_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_2,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_31: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"92225124929249248894408541300A6DB00792FFB12FE7240371F9F190FB007B",
            INIT_RAM_01 => X"0422500891088848884109240412044442091020842411042041088241144552",
            INIT_RAM_02 => X"9001624489A10045D16C944B02763FF55405E400BADFE5BFFFFFF00000000011",
            INIT_RAM_03 => X"49F30426B100842A12B25160D6D991E6C8C81AFB4C64400542140A342020D84C",
            INIT_RAM_04 => X"883838649E1442A3A1F70CA9094A5AD4A52D56C5D80CAC58D9645944A2300915",
            INIT_RAM_05 => X"A276585D5273AC87206840415DA74B4E9D213CAE3234B308E19608AA38250844",
            INIT_RAM_06 => X"B6E370363701B41848117683379C8422102D001BB41FB8248067301E1002C636",
            INIT_RAM_07 => X"84724A241226DB4809C9A1100DE6A63984D651A2624A09420496DDC12CC10964",
            INIT_RAM_08 => X"4C3C8D784218667F524CE209881213DC91099C14744901620044C802DA414966",
            INIT_RAM_09 => X"169808000200040100000002F8986E37654DDFF88E20860382DC089D4C239F6E",
            INIT_RAM_0A => X"1A55A50C3384B549B64C381920140D4008004020B119D4834C10064000006001",
            INIT_RAM_0B => X"0D1C3E528444D9B00E561C40973AE1806031C464834F03D34A11233A34B34A1D",
            INIT_RAM_0C => X"81E08228382D54C298DFC59535528176240438C9AA757917F95C7428981A2647",
            INIT_RAM_0D => X"184B56183004204267600220A061A004893E1D609106BDBB553920A011AA5AE5",
            INIT_RAM_0E => X"2DA65C2472B824F109BC594C2401209C01A0E59830002C73B396C6015B85A163",
            INIT_RAM_0F => X"101CC0024A6C32005CCB31908842211604D8B326101118B54B188CB4D502F5F0",
            INIT_RAM_10 => X"0BB04344008422327B1393C43396A931B8C8C87227A6141C0E2DCC76D830A082",
            INIT_RAM_11 => X"102B400E8004C40AD6E4614466308ABC7165AA57060A3A736A188ABB300200A1",
            INIT_RAM_12 => X"19B4C2CE666052C0619246C4B2245DE02B4009000402001E1051410804201E92",
            INIT_RAM_13 => X"000010004002001000200008000AEE708008880C86112252345B36C0048833B3",
            INIT_RAM_14 => X"0200080020000800200008000800400040002004000040002000020002000801",
            INIT_RAM_15 => X"CC0E00DAEC3000194A52B80C606262092D84A110241000000140001000200080",
            INIT_RAM_16 => X"10438134E31C28000400B18422CA60FC42C9C03F066366ECBBB010B00B004807",
            INIT_RAM_17 => X"881B30810845E6D18622EC9B6236A000030986A4F0644601226000A2F020C403",
            INIT_RAM_18 => X"C4C088B1A9B24BEB0178C4D6C18C3C5F72B07A28063647CC4721026D8C711864",
            INIT_RAM_19 => X"07D901787004001C459326210CCE00C6AF707B84440C313B10B8C4D13B2C6E06",
            INIT_RAM_1A => X"00800020249004081008924124080914000000020BFFFFEC638C31207B6C3214",
            INIT_RAM_1B => X"CB1E518948104042F84F1840401018402877D800A00000F5122597005DA44110",
            INIT_RAM_1C => X"6E436E644CF6C8D86F124DA26CE9B66E2F46BB466E2CE068661B4B05F02F7D00",
            INIT_RAM_1D => X"202139803D3000B2E0209DB9101160989A5916381001B0446631006064DB1B99",
            INIT_RAM_1E => X"C71478E35468600B01A93082C63DD073AE4181844449C08D8D56B0DCC881251C",
            INIT_RAM_1F => X"7C762E21DB2481CB6BB88C68811C76C63B18ECC1BACDC6110DCC70BC20940800",
            INIT_RAM_20 => X"66CB633B3376DC625DA8A0856C490392B779E1BA4088EDB4A6CDB9BD46DCC0B2",
            INIT_RAM_21 => X"FF7DCCEF40196C8381658D8840043B119B86A46247665810E2203000141023C3",
            INIT_RAM_22 => X"3124862592C0CD0F07A27A111CB80A48808C7C21C205029100010400228BB3BD",
            INIT_RAM_23 => X"C14D536A45D144B244C24A290076E58CC2E64E4A2DC4C5939C4C2DDBD1B918B2",
            INIT_RAM_24 => X"4B72C08871D2413188E4829219C38C2025920480D64856902E4D4D60B640C833",
            INIT_RAM_25 => X"2166D72DC524870C422BBFFD4808A7016B088DE3000B853800336C8E9968C19A",
            INIT_RAM_26 => X"C629E6050C619658692170C1022C2232C965C92C189020470587308485891032",
            INIT_RAM_27 => X"1B9CE2DA363196DC20007FF5554FC631286DC716B048384C26510685218DF9E6",
            INIT_RAM_28 => X"03C11245EE31E38E6DEF2188BE2068F3C716E10317783020D8EF5C256774BA0E",
            INIT_RAM_29 => X"7D8CDC0131C444798F040DC0116E2C4336B0166109A15D1FCC7EDE31EB238622",
            INIT_RAM_2A => X"4B987A78AE1BF80005EF370C0739371E0D3E5CF1E3677332370BB98D1831B30F",
            INIT_RAM_2B => X"0001022EC10015E263787F7E581EF83F062200C626EC4E19021840D9C112400C",
            INIT_RAM_2C => X"C23A8D170CED981891256A2C1D9B31C0F040202103900E6765976089DB8DE16E",
            INIT_RAM_2D => X"CFC3000F43632B49C39723270C604B184D1940F1B2A04459BEB088666943BB38",
            INIT_RAM_2E => X"AE6302C4BE6BA8C22A084803225A0855ABBBC528B1DD122B524A8D33C1209153",
            INIT_RAM_2F => X"873CB568FC3F09080F4400DAC600092017210911A6081DCC4979244124815884",
            INIT_RAM_30 => X"7FBBEC46E8B3CAEBE0100275A1092081D0C1E5716DF09CFEEC022D800529E1A8",
            INIT_RAM_31 => X"596CD8B4B568A4DFEF3DBF8027A3422A56A2C003E514582104BF8D6B5D80BB39",
            INIT_RAM_32 => X"0000000288964258156302504F5F660C054DEDCA20CC201A0206160601E376C9",
            INIT_RAM_33 => X"C7C57F084106FB3B8B1E47463C0088D11104F23C180222A0AA22A22882A202A0",
            INIT_RAM_34 => X"5775469089F04C623E19317B486F653C1C22CA642CD685C10EE47EDD66C8C226",
            INIT_RAM_35 => X"763C75FA1DB107B865E5B8F7B95E77F222244C6BDC1879C0562EF779BE000946",
            INIT_RAM_36 => X"06E5AD6C882882990A40D293FED064710CB226CDA0330D7B189B344442EC35E3",
            INIT_RAM_37 => X"03020CCE064769B15020A6030880234C64E9BEF8E98A81489083A026140D6489",
            INIT_RAM_38 => X"8C73E37081C37C37D6745354522D45157643E8840C02862C088C36E19CF1D315",
            INIT_RAM_39 => X"8C4902D2334D544B189717919B6BE6C731CC69288842152CD1857ED8D8E222D9",
            INIT_RAM_3A => X"8110200202D000093C44208838031005891217420084588B5F22850618945955",
            INIT_RAM_3B => X"800000006200CC62175193999098CB9324083858709866221FFC0FA000060103",
            INIT_RAM_3C => X"000000000000000000000000000054A0A65440E0748114449540F824CBAC2497",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"8000000000000200000000020000000000000000000000000000000000000000",
            INIT_RAM_3F => X"3C00000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_31_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    dff_inst_0: DFFE
        port map (
            Q => dff_q_0,
            D => ad(15),
            CLK => clk,
            CE => ce
        );

    dff_inst_1: DFFE
        port map (
            Q => dff_q_1,
            D => ad(14),
            CLK => clk,
            CE => ce
        );

    mux_inst_0: MUX2
        port map (
            O => mux_o_0,
            I0 => prom_inst_0_dout(0),
            I1 => prom_inst_1_dout(0),
            S0 => dff_q_1
        );

    mux_inst_1: MUX2
        port map (
            O => mux_o_1,
            I0 => prom_inst_2_dout(0),
            I1 => prom_inst_3_dout(0),
            S0 => dff_q_1
        );

    mux_inst_2: MUX2
        port map (
            O => dout(0),
            I0 => mux_o_0,
            I1 => mux_o_1,
            S0 => dff_q_0
        );

    mux_inst_3: MUX2
        port map (
            O => mux_o_3,
            I0 => prom_inst_4_dout(1),
            I1 => prom_inst_5_dout(1),
            S0 => dff_q_1
        );

    mux_inst_4: MUX2
        port map (
            O => mux_o_4,
            I0 => prom_inst_6_dout(1),
            I1 => prom_inst_7_dout(1),
            S0 => dff_q_1
        );

    mux_inst_5: MUX2
        port map (
            O => dout(1),
            I0 => mux_o_3,
            I1 => mux_o_4,
            S0 => dff_q_0
        );

    mux_inst_6: MUX2
        port map (
            O => mux_o_6,
            I0 => prom_inst_8_dout(2),
            I1 => prom_inst_9_dout(2),
            S0 => dff_q_1
        );

    mux_inst_7: MUX2
        port map (
            O => mux_o_7,
            I0 => prom_inst_10_dout(2),
            I1 => prom_inst_11_dout(2),
            S0 => dff_q_1
        );

    mux_inst_8: MUX2
        port map (
            O => dout(2),
            I0 => mux_o_6,
            I1 => mux_o_7,
            S0 => dff_q_0
        );

    mux_inst_9: MUX2
        port map (
            O => mux_o_9,
            I0 => prom_inst_12_dout(3),
            I1 => prom_inst_13_dout(3),
            S0 => dff_q_1
        );

    mux_inst_10: MUX2
        port map (
            O => mux_o_10,
            I0 => prom_inst_14_dout(3),
            I1 => prom_inst_15_dout(3),
            S0 => dff_q_1
        );

    mux_inst_11: MUX2
        port map (
            O => dout(3),
            I0 => mux_o_9,
            I1 => mux_o_10,
            S0 => dff_q_0
        );

    mux_inst_12: MUX2
        port map (
            O => mux_o_12,
            I0 => prom_inst_16_dout(4),
            I1 => prom_inst_17_dout(4),
            S0 => dff_q_1
        );

    mux_inst_13: MUX2
        port map (
            O => mux_o_13,
            I0 => prom_inst_18_dout(4),
            I1 => prom_inst_19_dout(4),
            S0 => dff_q_1
        );

    mux_inst_14: MUX2
        port map (
            O => dout(4),
            I0 => mux_o_12,
            I1 => mux_o_13,
            S0 => dff_q_0
        );

    mux_inst_15: MUX2
        port map (
            O => mux_o_15,
            I0 => prom_inst_20_dout(5),
            I1 => prom_inst_21_dout(5),
            S0 => dff_q_1
        );

    mux_inst_16: MUX2
        port map (
            O => mux_o_16,
            I0 => prom_inst_22_dout(5),
            I1 => prom_inst_23_dout(5),
            S0 => dff_q_1
        );

    mux_inst_17: MUX2
        port map (
            O => dout(5),
            I0 => mux_o_15,
            I1 => mux_o_16,
            S0 => dff_q_0
        );

    mux_inst_18: MUX2
        port map (
            O => mux_o_18,
            I0 => prom_inst_24_dout(6),
            I1 => prom_inst_25_dout(6),
            S0 => dff_q_1
        );

    mux_inst_19: MUX2
        port map (
            O => mux_o_19,
            I0 => prom_inst_26_dout(6),
            I1 => prom_inst_27_dout(6),
            S0 => dff_q_1
        );

    mux_inst_20: MUX2
        port map (
            O => dout(6),
            I0 => mux_o_18,
            I1 => mux_o_19,
            S0 => dff_q_0
        );

    mux_inst_21: MUX2
        port map (
            O => mux_o_21,
            I0 => prom_inst_28_dout(7),
            I1 => prom_inst_29_dout(7),
            S0 => dff_q_1
        );

    mux_inst_22: MUX2
        port map (
            O => mux_o_22,
            I0 => prom_inst_30_dout(7),
            I1 => prom_inst_31_dout(7),
            S0 => dff_q_1
        );

    mux_inst_23: MUX2
        port map (
            O => dout(7),
            I0 => mux_o_21,
            I1 => mux_o_22,
            S0 => dff_q_0
        );

end Behavioral; --Gowin_pROM
