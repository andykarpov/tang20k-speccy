--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.11 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Sat Jun 17 00:53:12 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(13 downto 0)
    );
end Gowin_pROM;

architecture Behavioral of Gowin_pROM is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    dout(2) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    dout(3) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    dout(4) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    dout(5) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    dout(6) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    dout(7) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FBE67965EC5F1297B17C565D9C5C25C3DD9F85C371AD97093F07050301A6EFD3",
            INIT_RAM_01 => X"7393118C96C0B703FC099189D52DF87E93342B864DCF5B29126DADD8FE3259BF",
            INIT_RAM_02 => X"F9FD7525CF0997298497D649F6DCE6597FD985C3D78AA098708888500AC219B0",
            INIT_RAM_03 => X"3AD9FEFA92A7EDBFFBF758CDB77BF677D5F7F8E522DB2DDFFDA93FFDF3CDD7E2",
            INIT_RAM_04 => X"16F95EE7ED49E7E99E5EA65DDFEBAF92689F7FB725C59277B72675573F8E522D",
            INIT_RAM_05 => X"2E9FFE007AFF4B328C0A77FECDDFBDF37EF6DFB35DBEC67DFBDDB3FEADBFC729",
            INIT_RAM_06 => X"07F7ECCBA707ABFE4927F993899F43FF99F4FFBDDE4D922647D68C279F77F9B8",
            INIT_RAM_07 => X"8A0CF9B3EBD1B6E712FFB23A5249F2192927D7E76633771FCC23A0BFAA798474",
            INIT_RAM_08 => X"3A03FBF6778F6BA707ABFE4927FA14BF987533EA7FE37FECE02596EAD8E2DB3E",
            INIT_RAM_09 => X"F46DB9C4BFC02A9E611D7FCD0342BE44D07BFDC7F3B31DBB8FE611D05FD13CC2",
            INIT_RAM_0A => X"1F18391FFA2A413166802AF764E64C0499A99E7966D5BAB624B6EFA2833E4CFA",
            INIT_RAM_0B => X"D2AB5AAABFAA8000039220C2A54C87FFE34BBA975B8971295BF897F10985FADC",
            INIT_RAM_0C => X"FC49624998A48F19629230402F56A9F892C70CC538714E24C31402F569BBB749",
            INIT_RAM_0D => X"446FEB2AC7081059B83D6558910044784C16F244E4C15A62532ADA4B0605528A",
            INIT_RAM_0E => X"7FFECC6F3BCEF1AC6338CE779DEA715A7370F918A60371ED4841B9BBA9082E5E",
            INIT_RAM_0F => X"00AFFF4040A1F7BDE615A884831196498912510FFB9FFF8DFFC7FFE37FFCDFFC",
            INIT_RAM_10 => X"0C37BBCE6A4C4C4C7D95537AA64A4E54F528532DE261F7FE682187BDEF320F02",
            INIT_RAM_11 => X"E3CEE39A29C6B1E13CDCA9352852AD5A002AEAAE615A8A26AADE48008495FC11",
            INIT_RAM_12 => X"149B3AADE970D909DE72C9DD93B6D31E9CFF2F3601E1BD494E6BBBF9F5DDFCEE",
            INIT_RAM_13 => X"D5B9EE0DA473EF60C1F9B0645B77ED9CD505C8CD2DF647CFB31DBAF58D84067C",
            INIT_RAM_14 => X"AD8987531E9BD9D2EFFDBB7B7F98650E987EB7A7BB66D576FFFEA4D275082E1D",
            INIT_RAM_15 => X"A4B7AC94490D59FA0927CF22C54CE299E2E01AD7DEDF5D5BAF234D37FF7FE6EB",
            INIT_RAM_16 => X"DB8505264C0962D2EDDAA668C982600A8281748C0D73AEC860C08AB6056A18E3",
            INIT_RAM_17 => X"F276C12439CAFFF7F22AEE9144511114077D82C987A091756A272C11C208E5A9",
            INIT_RAM_18 => X"7FBCC602B477B3D9ECF67B3DBD3CCEED092DF5B56967584DA59FFFF75FA695C8",
            INIT_RAM_19 => X"40374FBFE73D1B0BDD277C4E00CFE933560F6FEFCE4E62DB39E1695B9EE1BB1C",
            INIT_RAM_1A => X"406208040241248049041041046A371D700001B9BA4DBBA613999AF6E5DB8592",
            INIT_RAM_1B => X"52D4725AD5BAB57A24AB528DAFF86F56B5AA94A52E9D56010124043577616400",
            INIT_RAM_1C => X"E9D5CA75729D5FE7C93F819D46E33127485B81129083EB850165A4346A5C04E1",
            INIT_RAM_1D => X"036A4280882664D4D4CED9A7CFF11DBA74BA498A7263F9159FF3C9F7EB679F27",
            INIT_RAM_1E => X"F9F9A4A4A4F6BB6EB076349F3EECD9367DA4D6CDFE1C752B29997961302B1B50",
            INIT_RAM_1F => X"FBA79847407F7FC91E0E33E4783CFF353B3000EFCC25862402D95E0004C25809",
            INIT_RAM_20 => X"516014F092D7C32ABDF9670674AE745C5C966593940824BE4FF23671FCC23A0B",
            INIT_RAM_21 => X"963B9BEA7FD5B0A4402D4A2B659F3371FBFFE557D9739901264989FFF3C0C0AA",
            INIT_RAM_22 => X"D365E68B4D8FF2C2120F49C83D3722FCDD8BF3610D332274CC89D13607C4D83E",
            INIT_RAM_23 => X"5D7FFF4D29345A6858DD4BD18CD33ABE9B6DB5643EFFBE1CF2DA1B3A5E5E94A0",
            INIT_RAM_24 => X"B52B339FEC98757379316BA0665E4F262717DE7F5C077CF2F34F673ED8FF79FF",
            INIT_RAM_25 => X"4E24D3FFC1BDF9BB344842E75DABFF778FD99B326A8B9A482E6908A0885D4150",
            INIT_RAM_26 => X"FF1924386D059751F70F309F85AB818CEC800099966671989BA42D00C0B5C652",
            INIT_RAM_27 => X"5AA4A12A4A132923773EC1D0D9056FCB8869E19E87E79CC754CD80AE669F85E7",
            INIT_RAM_28 => X"FC7A2EFE5FFA7F16A6BB43B3308EBCED4F3B53DDC73F36D4F307CDA840040110",
            INIT_RAM_29 => X"A802A42C054448192A2028C4883C38FFA7DFE55404BE7D76D95A0112ADF7D361",
            INIT_RAM_2A => X"06A4894F84B955670962B639F34B3E717AD230A77D6CE4EB3CB1C76F18702A80",
            INIT_RAM_2B => X"BB5D1976CFFAB6FDF1339B21375D81FF649F1CF8927DDDFCB36EDD3C9D044C8D",
            INIT_RAM_2C => X"E79D36F7ECE7AC8B74EFFCD1B3FA35C69BB9E599BACE6D9722D9937AA99263CD",
            INIT_RAM_2D => X"FA6CDA265930E691B3689964C3EAD9BA3C003FB96887CC5BAFF3474FE8DF1A6E",
            INIT_RAM_2E => X"323BCC5BB77A4AA5162960C8A12DAB6CD9C6936D99CD9A9F349C921239F8B3E5",
            INIT_RAM_2F => X"1C1C6F0F3BAEF9ECA70EB7E726F61BD21FD21FDFDDD66B09DFAECC14879FCFCA",
            INIT_RAM_30 => X"2FD666A9DA26BCC431766B6165BF26DB3B70923B7FECA1802EEA8BAFF4FAC9F3",
            INIT_RAM_31 => X"33326E9B6D94291EBD864C9BA7723A2D47A49F5219CEEEC1204427F26D2166F0",
            INIT_RAM_32 => X"B86414C656787F74D27C6984031FC5B369D253CE9CCCED0112042CDE77AF3333",
            INIT_RAM_33 => X"4B5B6A080D38A040C8A42E1E12832BA2134B5CD33A490DA5AB3A095522C0F375",
            INIT_RAM_34 => X"1038B2A9D136825D3A3A1B0C42C924752AD0A904A85540955055B06218C562BF",
            INIT_RAM_35 => X"33285A224A25932CD01368023C584003C268954084AA18049371A408345080B4",
            INIT_RAM_36 => X"849356CBDF4139AA08AAAAAAAAA00028225FD75F57F7F77F7555D6A2A8AAC2F0",
            INIT_RAM_37 => X"71AD6F7A539353A4B7FA27D614FA46751DA4D26B5CCAF892AF2B2A4DB7BA9D78",
            INIT_RAM_38 => X"0244441DFA9BBBC2222266CB9ABDE66CB99BE1062538E6259CC9B76DC91DE326",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000001400000000000",
            INIT_RAM_3A => X"FE00000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"0BFC000000000000000000000000000000000000000000000000000000000003",
            INIT_RAM_3C => X"87B1A2222220F8687B1A3622220B8687BFA3622220A8683BFA22220882838FA0",
            INIT_RAM_3D => X"000000000050108A29A0222210828888888200A22362203068700A2236220FC6",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"E900000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"12A015843641BB14D946E041A2C10C114242240267194B027301010100538761",
            INIT_RAM_01 => X"AC4222620115A15D41C4AB0F9EFA074004573E140A163A9004F1300FC3073034",
            INIT_RAM_02 => X"2E42592E2EAE1CEE381C676E5CE3B0A1C25E2E10478FE14AB02829140363653C",
            INIT_RAM_03 => X"0CE7600398C61E7BB7CB2F163175CDB195C170E62198CE7602399623CB8E761C",
            INIT_RAM_04 => X"0CA643A011CCA1125C43A1834212CC9616A5D774A2A02A1754DA1954170E6219",
            INIT_RAM_05 => X"9005D1AC480721F039528D410A1CEA2871A0B544BA5578814BAA6D4CAA0B8731",
            INIT_RAM_06 => X"A2201921562B5200900818ABAD39ABFE9E6F35401AA254641A043F1725C0AE45",
            INIT_RAM_07 => X"4AA20A9224A29206889B16683490C1501A4B3840C21D645196CD75D11C32D9AE",
            INIT_RAM_08 => X"D751100CD4F0E1162B120090081EBDD98871A7317FD34C60ED03CC40C56020E4",
            INIT_RAM_09 => X"28A481A23FA052A4B66BCD9522D641A0B5652A7A206102B228CB66BAE886196C",
            INIT_RAM_0A => X"9C8340BFFAA8D7C398F04C5C50B45365A2922B04404310314009B912AE82B489",
            INIT_RAM_0B => X"FC675CC67FCC8000020973E7EFFFA7FFEFF8988E183B07441803F007C0A9C6E3",
            INIT_RAM_0C => X"C01E1409A5E8065017A03F0018649D803C2B4D2E580B9609C3F0018648E37867",
            INIT_RAM_0D => X"6C4BA0A22B04C97128341445008E8A1C75D1840960281014184C811850833646",
            INIT_RAM_0E => X"62AA028252842319C63084212945E19262560305DAE25758F21129311E4424D4",
            INIT_RAM_0F => X"64202216742A27C60CDFB116E630496C459463517C1CAA8E55462AA31550E554",
            INIT_RAM_10 => X"D557CC180779EDEDC60642C0FE8F1144019B340C16081810C33B293E3067BB64",
            INIT_RAM_11 => X"9B32C731260FE06B7C2288419B36895D21B8B7D0EDFB12B6C810DE4116C40129",
            INIT_RAM_12 => X"5D4843FFD3C4549EA4C3D1921F330B3921C806987B54C444DCB7FFFB1BFFFD8B",
            INIT_RAM_13 => X"E724409CD38A088C2CF2BB268B152E204476AD4DAE446A04A17529A05E20C4B7",
            INIT_RAM_14 => X"009A23815508561D00C44E0AC4D192105143AD02A4A14852843C2852B50FA8FE",
            INIT_RAM_15 => X"32286884324650726072786B41FD43FAA06B2800400120442A73C2502ABC0FC7",
            INIT_RAM_16 => X"92264064C11010166059850E459A12D88680AC55990348800402BC1300402920",
            INIT_RAM_17 => X"01355069701189EC9E3AFFFABEAFAFAEF3B0CBD9D609CF1D7A4E48B002180509",
            INIT_RAM_18 => X"F92019B371E4321B0D864321BEC002DAC31BA398E64A3CD28C08860C06E7E8FA",
            INIT_RAM_19 => X"C012013FEA51A4C760D032CF547D4683554034341C002607564306308FCCA098",
            INIT_RAM_1A => X"41640904820100020800120120C25984680000E00320E080A2AAA519B27648E4",
            INIT_RAM_1B => X"64B028C28428A4D2194840158B31456739C98C63008953402000886165A16092",
            INIT_RAM_1C => X"0A2412194CA2434286D403003D100BC2210808500999C8886C41144C266B042E",
            INIT_RAM_1D => X"9A2D875E0B04154B535266E0212BC854A810F298BCAC9B37349614A4321D0A04",
            INIT_RAM_1E => X"D1528000000970C64D8D900C18964E1E207863C626A075B2283831403180916B",
            INIT_RAM_1F => X"11C32D9AEA2200911E5D9D847972447C7832E5E6001400A0C13B610CC08406C8",
            INIT_RAM_20 => X"C8E03A023C2F68131410A0FA0EA89E40581C110054B9622E0030D745196CD75D",
            INIT_RAM_21 => X"8E5F12EFFC41D362C5919063815468D4054C0262A2A2D0D9688DC149550A1066",
            INIT_RAM_22 => X"C1B78B6F84C6C0010675C6B8D30E61C4B8975020032AE55C298730E61CC7B89D",
            INIT_RAM_23 => X"14A1874B090592496AE18C18886F69990C37D97C43237DC06F488008E1872DD9",
            INIT_RAM_24 => X"19A547A089A2381FFA020514AEC2DF5A066E0003FFDFFD37F4908F45C5485844",
            INIT_RAM_25 => X"9C09E841C8494B18D727266EB0954604D92BE1180545B68A16DA204049E8A351",
            INIT_RAM_26 => X"1350D1406D08DE717556516F952603BE03AD6FB401D38C05CF1013B9858D80D0",
            INIT_RAM_27 => X"4C5294AF6BDAB5A99FBC3329D89C8FFE30002ABF3800B3FAE605D41B00C83A01",
            INIT_RAM_28 => X"06A12CC0401F4982B7815BDA5B35D0056F815B80016082DC003820A456B5ED39",
            INIT_RAM_29 => X"3210CD08C068B20A8808002804647400B0001AAAABC8F7E30C133C10D8C22608",
            INIT_RAM_2A => X"0EDA0514C0DF056181A95CEE2A2F7B19CA5074FF1E999815888AC75090040B41",
            INIT_RAM_2B => X"6B2EE2B1B632B02E41BC8C0171DE65CB181CBC410B61E361431C50A06188C827",
            INIT_RAM_2C => X"C10AA25442A10A91205552E395790C2F0EF041A750AA1014102A6D4CAA020341",
            INIT_RAM_2D => X"1933C5FEFBFDC33C4F37FBEFF7132F461460AD84F1E80E89014B8F55E434BC3B",
            INIT_RAM_2E => X"E9C702D28151066C8E1E1AC6213FADC32E88FAA44E895816A505B6BCEE295C99",
            INIT_RAM_2F => X"3240B15CC109C58AF79F91A90A3A7DB679B679BEE95EC3C1CE0382A3702DDB00",
            INIT_RAM_30 => X"A5C69A8ECB72F9EF4AB02E434C28D3C0F08D81209912E3871A115F989C0150C1",
            INIT_RAM_31 => X"41410BD1281D7B87EA74042A1F09069FD51A592AEA1B48222CD7B4CCBAC4430C",
            INIT_RAM_32 => X"38B01FBCC3157D238E958C2D5604E89A0E3380918525148825AD600520694141",
            INIT_RAM_33 => X"2A925198DDB2306D06664CA1A78A33121A5A8DB32215092D4233424D91A08846",
            INIT_RAM_34 => X"0940A808593E91514328D1C4228A2E5848D3B6C6AC028B80A10524A7086762BF",
            INIT_RAM_35 => X"A098C6444C6106188C13D818347C10084F380C906464831424336D845A310020",
            INIT_RAM_36 => X"4D3FECADBA07C52AA82222228A22000A827D7D7F7D77DF57DFFD5D7557403060",
            INIT_RAM_37 => X"88B1B476B5A025CF0803FA8A62156CF12C5A8AB27678546452B17801051384B4",
            INIT_RAM_38 => X"029414F32D92C1957D7C29D96E8B029D96A99456E85644499B93E20ED0C482D5",
            INIT_RAM_39 => X"7010604000000070D018C0C040D13000600800200000000000008088C0900000",
            INIT_RAM_3A => X"FE0020010001080189F838F800C1117030F1F9F90100F909F9E009086090D1E0",
            INIT_RAM_3B => X"0BF80800010801F110F030F0808003F060E1E1E00001E801C1F00121F8A0C1E1",
            INIT_RAM_3C => X"0FF900000003FE40FF901400003F640FFF81400003FE40FEF800003DE00BEF80",
            INIT_RAM_3D => X"00000000005037A69A7C000035620000000DD980014003BA409F900014003BA4",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0C80000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"4482A1A97685BAA5DA16E2050E050151072721448460879FE402000200D691F0",
            INIT_RAM_01 => X"E8893344D015C3D10755AA229E322684099285341290A9093FDA3555471740D1",
            INIT_RAM_02 => X"A2A9A62956B28572F205DA62EE8583001752E150C0A1441AC002A945000F40F8",
            INIT_RAM_03 => X"9F0B04435CE172AEF61492A2C35C1C839615D846116572F15635F1561582B97D",
            INIT_RAM_04 => X"8B6BA792B1AF92BEAC25D3B7254D3195B34EFDED517349B5CD89B16D1D846116",
            INIT_RAM_05 => X"368F76AC58AF6BDAF15D3C9106E166AD8792A4D536AC95269AE6E49CB6AEC230",
            INIT_RAM_06 => X"A2A80B42E92F41FEDC18B8B484FBB4FE86EB726E79B502221882B6058C9D26ED",
            INIT_RAM_07 => X"DCA9B3C49B3BD3488B3B1069A490D814D24BFA810212122C0CABC5D55A419578",
            INIT_RAM_08 => X"BC515405C5D482A92F01FED818BCB9FB80909F709FC01CE009024DAB90F72AEE",
            INIT_RAM_09 => X"CEF4D222DF608A08655E1DA83496C461257D62EA40810109160655E2EAA520CA",
            INIT_RAM_0A => X"D7AB008007B216E0CA5C7C4518535FF508B088A822036AE425CA1BB7286CC126",
            INIT_RAM_0B => X"DC1F5F01FFF0800002031364589025554D91830B61B636C5695B32B6402E1F0E",
            INIT_RAM_0C => X"028942409004C22D40120FC20F6BAC051287C4823E208F7F80FC60F6B9A6EFDB",
            INIT_RAM_0D => X"E0A43C8087B0B68290079010960056E8F000F258F3A0EF425B961D40A100F110",
            INIT_RAM_0E => X"A6AAE6E842000000042000000006038805202374D2052460498292440930D04D",
            INIT_RAM_0F => X"4520221494EA27C40CDAB99A45304A6C95F67B517CADAAD6D56B6AB5B5554D56",
            INIT_RAM_10 => X"5D57C81A0B8870714600924AFA8F53183693252950A85810C24B293E20671C45",
            INIT_RAM_11 => X"D29EA61A139C382B7E1A3056932E440F31147D5AEDAB1884C30EDC4116C40122",
            INIT_RAM_12 => X"DF6E83F698146082B6E3949BD9274A31B52862B86035C1859EB000029800015A",
            INIT_RAM_13 => X"58E82A89CD3E87882BD21A0ECCB432A154224DA1B2B36C40C53F09F142A05285",
            INIT_RAM_14 => X"2C06A3E14E2854DD8AE56CB8DF4CF38DCD3D8D8126EB1510DFBEA492791760A5",
            INIT_RAM_15 => X"EC12A184AE1E01892536E04B6DF56BEAA64A22D51E94540B6518DB7A1141B2BA",
            INIT_RAM_16 => X"992204044990344440990264D8B1608234C2A6C404A1C21941A13D6903BE4243",
            INIT_RAM_17 => X"7845D875705A1DE9D62AAAAFFEAAFFABF38580495262EA366A0EEC89A244D084",
            INIT_RAM_18 => X"81B45F3875AE030180C0607036AA8237470975394E2750D10E09CF204620EC33",
            INIT_RAM_19 => X"C014448AAD6DB5C2576774A45475FB35FD4149497C00057C7B22BB508F29BA0C",
            INIT_RAM_1A => X"00064004900104104800124800349288100001A5BECDA5B6A1BBBC5428400A86",
            INIT_RAM_1B => X"6954D21975C65D6A572D5F0F2E58BB5294A5294A14D0000903248C1A09400482",
            INIT_RAM_1C => X"76FB7DAE974BA7CB81BEA8EC767D1B83583B6112B28131160FA48874AF61168E",
            INIT_RAM_1D => X"1DC4411F852B405CC4C7298F53B267783842E0167A69C22EA9C793FB7DBF2E03",
            INIT_RAM_1E => X"A0022020204DCEBE55AEA00C5C1F0F1EA7FC7FD6762464333890C0B6581CAE20",
            INIT_RAM_1F => X"552419578A2A8118A69D8DA29A72041C194489264464872401C326001614E408",
            INIT_RAM_20 => X"22000809128BAA3F117083E8BEB2AE04502000805922401E0170A122C0CABC5D",
            INIT_RAM_21 => X"1000296FA159E74F9F9CB112C3D10A40535143E20AA94DF94206C21C4554201E",
            INIT_RAM_22 => X"80F749EE1143A041180E01C0380300608C11C2008C0780F01C0180300604C084",
            INIT_RAM_23 => X"4496F7631915D96C620A730A101C9205830FC57A4777528414C38812AF8C0B79",
            INIT_RAM_24 => X"78234736E84A3E56D3C964EEE0AAFA78404E275AAB8AD5B5A6DBAE7E2D37788F",
            INIT_RAM_25 => X"FA7FB8E6009494FA878D857CC42359A3D1EF3E1C2A9050024140090901E2A040",
            INIT_RAM_26 => X"3AA02C487C5E555D459C78E292EB0329AE3ED28C856D3C8DCDAD97B124152667",
            INIT_RAM_27 => X"1C300C010250A50B9828A299148A6ACC9688EABF2B62BA60D480D42B02E3A861",
            INIT_RAM_28 => X"7E8B2C90856D5DD6291B102432AF166C539B140DC20D96003193458610806018",
            INIT_RAM_29 => X"120C4CC6C6CD731E20A0A084B4090B02C38B40000140EE471DEE3F0A40C630A8",
            INIT_RAM_2A => X"0ADC993D44F3657C89F17112F9D548A8185666FA2D90A8375C21EF252CA42100",
            INIT_RAM_2B => X"401254839172C2A2A14101B94212B618B205582CE3050F0600B7DD4C07244421",
            INIT_RAM_2C => X"E00C974D8253AE6BB1741CE841A01B400FF8014BDAE9B00D39A6C498B681A335",
            INIT_RAM_2D => X"A84B53CCCB7DC6A9AD4F332DF74022DA1620AAD1B52CA65D8873A006806D003F",
            INIT_RAM_2E => X"B69F46E0C19AC1E220094B82E0AAC28A6EED38F54ED1048AB98DB4B916F17DC5",
            INIT_RAM_2F => X"2860935A2F894EEA159B9421128861646564656DAF1A019B452280B0CA8FC742",
            INIT_RAM_30 => X"248028041BC05DED5D54A880013E2E02D2DDE532BD12020112328FA9DD3AC6E8",
            INIT_RAM_31 => X"111859EA3119738E12A8044BBB59ACDE9785EC50019FECF2ECD538B01E2041D6",
            INIT_RAM_32 => X"82E77E7385B29D5716A01D0957A0351DF2F140D044544528152D613074111111",
            INIT_RAM_33 => X"81C832085096910E4AF6C1269A85B6D00839428384D0041CA20C8D20B4224C37",
            INIT_RAM_34 => X"08489169DD38C2451018584630C3267D92A33740AD3AE34EB8648CA321E13417",
            INIT_RAM_35 => X"59A80AC09C6E96A2EC13A81979C5700160081A01A6D01D15A1050550E00429DF",
            INIT_RAM_36 => X"94D7BD54ED213A822A8282802A00880A20F7FDD555DF5FDF5DDDDD5DDDE72184",
            INIT_RAM_37 => X"E78289100006DF64A7FF242B5D460C40783CE8358CCD829D3D35CB3EF86FC889",
            INIT_RAM_38 => X"022BFE444FE916157FD4AE1B0F31EAE1B0FB1C7300C22B9AC1BF6D79E9E5316B",
            INIT_RAM_39 => X"7838F040000000F9F839E9E9F9F97900F01800200020A0600011D159E9F83800",
            INIT_RAM_3A => X"FE00300181091819D9F879F809E9B8F879F9F9F90189F909F9E80908F199F9F1",
            INIT_RAM_3B => X"0BF01860019913F1B1F071F101D013F0F1F1F1F10113E801E3F00971F9B1E1F0",
            INIT_RAM_3C => X"16AD060606079301EED074606069B41EED834606041B01EED8606040101EED80",
            INIT_RAM_3D => X"00000000004577AEFBFC60604010181818140406034607BB4168506074607BB4",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"FB00000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"408A81E862948AA18A522A9508950951066F294190C411C26C000200014624D0",
            INIT_RAM_01 => X"62E1113490B38365079591E27C11A294499784C912C4282084D56F761C30F090",
            INIT_RAM_02 => X"B282DA5856108560A3212880A29683821F508951CF605A56D0000051402CB0CA",
            INIT_RAM_03 => X"142B044B9EE852A7725C202242EC188A2C58AFBD2C8142B044B9B9421580B151",
            INIT_RAM_04 => X"640A058A25CDC218AC1582338416D52C2D2A2AA1820320AEC58822C18AFBD2C8",
            INIT_RAM_05 => X"5E9BB98FF2FA485211C0AC5112856288158A24D112E101021760C45162C57DE9",
            INIT_RAM_06 => X"21FF80D087670600C806E8433C9B830EE2E9F328F9940E42058EB18EBC5122A9",
            INIT_RAM_07 => X"0C509153C911DB6D0179B2C362585A01B12F8BA323AB66610E2AD1CFEB21C55A",
            INIT_RAM_08 => X"AD10FFC04D6990EF676600CC06FE1CAE8CE79376E1CC9DA22C024E1090319E5C",
            INIT_RAM_09 => X"4476DF405EE112187156FCC96F873743E1F366B4D191D9B330871568E7F990E2",
            INIT_RAM_0A => X"2BA718307C674A4DD36E7A4952468A52EE5EA9BCC243842400671703162465F2",
            INIT_RAM_0B => X"3757FAB57F548000038371624C9E82AAA57D398A3B13624733F127E246C8966A",
            INIT_RAM_0C => X"C0084001B0800A41420130442D30298010818D840C610309A30402D3018B6CC2",
            INIT_RAM_0D => X"C001A60C81B024880034C190060E200871D2D008350800401A84445840A00480",
            INIT_RAM_0E => X"A556EEE10852908421094A10842A95011006032170C000C4400000CC88005240",
            INIT_RAM_0F => X"26DFFFCA1B45F73AE6F23DC8FC388E37DC53582FF3A95594AACA55652ABD4AAC",
            INIT_RAM_10 => X"60B735CE21D97839D985D2D0EE7ED64C739327A844A8E7FE7D0C97B9D730784F",
            INIT_RAM_11 => X"D18B5BDC712614883D3498B3932507799D58666047235DD99008A87D5B7BFCC8",
            INIT_RAM_12 => X"EA265FBE8A5622101A32CC4CA51F2D9CBC6F4CEBB9C3DCC18E8AAAA9455554BE",
            INIT_RAM_13 => X"4C8E7117CD2884044BE0812C08B1A2F1323B4D9A62AE6E460088045B12A0E2DC",
            INIT_RAM_14 => X"8ED0A2A4D82200653200241046DAE3A49C6D044002402D4A546880401C1E3784",
            INIT_RAM_15 => X"60042616A3428524496DF34681DC87B9D0E2B891CCC718E2D5D2E96B19BCE09A",
            INIT_RAM_16 => X"DBB563668C0B103668C0B56A15281051B2D2D4D9123872606400364804010042",
            INIT_RAM_17 => X"21459D9930D7BC07C20455111044441106CDA81840B8AB36388C4902D8816D6D",
            INIT_RAM_18 => X"D09E4B555F6379ACDE6B379AFA6EC024A21118FA3EB450C90B07DF6C5430A080",
            INIT_RAM_19 => X"FBA64100116BB96283B57D6136179DA4A9277B7A7C260F354DA79D54414D1354",
            INIT_RAM_1A => X"0904492000012080000480000080151400000189A60D8B3171111B6D9B369E60",
            INIT_RAM_1B => X"300000501514047351CE41074AA1124E739E318C288041810304044053800480",
            INIT_RAM_1C => X"66B259AC966B2681017AF4EEC65D028059098C40809B82C26C082141463406EF",
            INIT_RAM_1D => X"188C87008200462CECAD39CE679E63209947323C7E6FD37EABD5837259AA040A",
            INIT_RAM_1E => X"3C00A2222224D38E77EC3004488B251E215425C6F43657BBA018000671860463",
            INIT_RAM_1F => X"FFB21C55A21FF82D18BD0DA462F0045E59758B26C5049124C103340CC86232C8",
            INIT_RAM_20 => X"906038021080A0BE116082C829662C97E4223301C962C26607DA377610E2AD1C",
            INIT_RAM_21 => X"D69C801EF111B4A85049F82362B3A20A1B8873D209891A94BAAE225641481400",
            INIT_RAM_22 => X"24DE01FC038320A2920E41C8392324740E819051490720E41E81D1322640C82C",
            INIT_RAM_23 => X"52358D47B97492497BAC63CCAC11A6840309A78B2E71520C18A701060509296D",
            INIT_RAM_24 => X"0A8B52B3A12A2A022B1071A6CAC845695174839215A62D90565E2566086B3009",
            INIT_RAM_25 => X"9809A3ED08181A300EB6AF23325384A208488300044ED3243B4C90D0D1B68071",
            INIT_RAM_26 => X"7BB82C6C7D8B5555554514620023D18989EBBDCAEE6D2A81052D9FB1C4A1C090",
            INIT_RAM_27 => X"DD5AD6F5AF7EF7AAB55EA3FDBBDFF7AB9C08059CC9E38C42BCC4862890612422",
            INIT_RAM_28 => X"2261DD9AA6BEFC654EF2B7B438AB75CA9DF2A7397267854C7139C15F5BD7BDEF",
            INIT_RAM_29 => X"1B00680080481A1A202020803854406A90C9B555547A5D1DF5020100CECE15A8",
            INIT_RAM_2A => X"0E78C1110297193A052529E4F4F559BA9CE476EFE2F3A4529C20660800442B02",
            INIT_RAM_2B => X"4924049B134593348FD30952D314D2D92329E06D7435493705B4C9446F1C8406",
            INIT_RAM_2C => X"A3864749C09A25639823EDFF6CDF1B7C8DE8E16C8279302941A4C4D166C53F24",
            INIT_RAM_2D => X"EA4F5BC2DC58D4B1BD4F0B7163461DD21400ABB98C9EE19CC3B7EDB37C69B237",
            INIT_RAM_2E => X"369740800042C00906084384A02AA4C306399470463CFE0A958C22A9E6F52DE4",
            INIT_RAM_2F => X"EB5340703642CCA2758B0408480931E435EC35EF211CC79787A18688A22FE777",
            INIT_RAM_30 => X"8E4EB99A90A2B0755A40908209122E46561E05967C827983080253F9C1319000",
            INIT_RAM_31 => X"9994E8C2001C390A62AE00213A150D43B245C5126807259FC2AD1CC89224B500",
            INIT_RAM_32 => X"52DBBCC7052AED073833BD1F350E2908C2A4A4078A4645380DEF4044C1AA9190",
            INIT_RAM_33 => X"E08004008004000C2266493482081A20E01856999018700C25A00A1422C0683A",
            INIT_RAM_34 => X"006C802A951A994D089259800000249880831E0288670319C0184A4634402005",
            INIT_RAM_35 => X"81085048E86027049051881BB9C48009C330D55406AAC4043055240240563400",
            INIT_RAM_36 => X"0415EE06EC4D1017DF57FD5777D75F7D7F288A082200A2A28A8A0088A0818000",
            INIT_RAM_37 => X"22CAC41318CA054427FBA16A40880E46290095180CCA200614198D5422429580",
            INIT_RAM_38 => X"024444089D800017D5554818062DB481802B534A3269900891D3708860D01400",
            INIT_RAM_39 => X"697998410800A1A928692929F9294901183180208020E0F10819F8B129F819B8",
            INIT_RAM_3A => X"7E0019F8C109383870C0E1000928E9C84908E03101D901F82128292999092859",
            INIT_RAM_3B => X"0BE010F1F8F13280E100C101215010909110101101B200002290295121112150",
            INIT_RAM_3C => X"1EFD86060607FFE1EFD874606077FE1FFF87460607BF61FFF860606BE61FEFA0",
            INIT_RAM_3D => X"000000000048928A28AA60604A8618181812A186074607FFE1EE986074607FFE",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"9800000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"520A80D06F179141AC5A038709161040040B384446318A008706060401B10023",
            INIT_RAM_01 => X"D2CD33A6E49D0A800404897E1C7170851987F48972D0B317010A0AAA8824B000",
            INIT_RAM_02 => X"128187207712E140A165585085940A861B32D040D83C4E02C2AAA814503126A8",
            INIT_RAM_03 => X"1128142B9CF950E0BA50C201425258430258174D14A5108042B9A8421DF2A050",
            INIT_RAM_04 => X"A528940215CD4A10EF950A02840C359029284121442030252584B0218174D14A",
            INIT_RAM_05 => X"44794A855EA8386E1F04A010B2A50084940A10949286101A1292C21812C0BA68",
            INIT_RAM_06 => X"07FF385AA8670C004838A054CD9B84F602ED41086014742464DA5C15085400A8",
            INIT_RAM_07 => X"8C21B345DB33FB688BB868D7824857ABC1250AA121E1F76C36CD90FFE8C6D9B2",
            INIT_RAM_08 => X"D903FF9C05209AA8670C004838BBB6E20E99B3729EC05C838E2341900540086A",
            INIT_RAM_09 => X"CCFEDA22FDE20AA9B66C9C2664001539002140905090F0FBB61B66C87FF4636C",
            INIT_RAM_0A => X"4424482000C052224A426C0109529B68C85C802DA45064015C029AA3086CC176",
            INIT_RAM_0B => X"E0CFFCCCFF988000028159B068D4B80006E54B0C69BB37C7695BB2B7C082500B",
            INIT_RAM_0C => X"009615C0246B857411AE003C300D08012C2A01235008D4020013C300D0408235",
            INIT_RAM_0D => X"229E20302A00DB627804060570009C06800305C146882415C21A894850EFF700",
            INIT_RAM_0E => X"06A8E0EC6318C631842108C63185E6C644F030510A04F630B2027A221640A891",
            INIT_RAM_0F => X"06A81FCFB0E5F83F02A237C054288A64E847522E82C5AA20D5116A8835462D51",
            INIT_RAM_10 => X"C4B83E023BBA7675DB09AACEEC2E93D826DBBD3A49A06C0E7FD997C1F818500E",
            INIT_RAM_11 => X"93A0E3F474476420FDEBB006DBBD128885912578CE23D4883A64C17B564500EE",
            INIT_RAM_12 => X"0F0E1BBB64D060E440DAC6B014092B589D23D89AAE845584E25C4403AE2201D1",
            INIT_RAM_13 => X"9A489002518CB2D42C20C93641A484E027234D9046BA6D42C417209C26C2E94A",
            INIT_RAM_14 => X"6466C1E12F08443C098468188929E7FFA8B18DC209225259D0420BD0A518DD2D",
            INIT_RAM_15 => X"1A2B499A140010C0054B39F665D863B030E48F4C7239E5AC5552993A6E80B1A6",
            INIT_RAM_16 => X"8B366424481130444C89366C99336482A65008C8189A009067C3812000902325",
            INIT_RAM_17 => X"2438AA08319DADE6D22AEEBEBFAFAFEBE230410DB419014C62E099EA22F51D89",
            INIT_RAM_18 => X"C5BE5D7169672B85CAE570B878484B1221134C5B16D935BE1602D35C86DDB412",
            INIT_RAM_19 => X"731080CAA16DBD26FC9A2A77263B24DD55265A5A5E2E27CF6483E495CFEE68EC",
            INIT_RAM_1A => X"095800000238049209E4924927F644106C00004011A0419C0D33325123445CC0",
            INIT_RAM_1B => X"0DA3ADC7A079E8850A108C581187843DEF78000016431830E0E303FB0E1F6002",
            INIT_RAM_1C => X"76BB5D2E976BB5C3047FB64909190BC130306B10BB413A1800995E08A10A78E0",
            INIT_RAM_1D => X"04208400723D13AA226134D2658F649C3849701E9A8ADA3F36D7041A5DAF0C1A",
            INIT_RAM_1E => X"F6A84040401270C14588508C182706202058C104B083AB5547E835D000002100",
            INIT_RAM_1F => X"FF8C6D9B207FF384A4BD0F0292F00E5C4845AB6EC411820C002841001A900202",
            INIT_RAM_20 => X"E00020032C2B029B01604A442416A185542216829962C2DA0DCE1E66C36CD90F",
            INIT_RAM_21 => X"1AE627AEC9C2393264E8C804606228085801776008054ADA322E641A014A1DFE",
            INIT_RAM_22 => X"80A301460040A0411E6FCDF9BF33E67CCF99F3208F37E6FCDF99F13E27C4F891",
            INIT_RAM_23 => X"9656082064410925AFAAB54C05A690480453A94F0AB1E56421308F30850D0D53",
            INIT_RAM_24 => X"002000724A2C1E5807432287EAC600F91C67234C108407A00E4EACE940B4E809",
            INIT_RAM_25 => X"20021165081A5A0A028E27C26A4010392D409130004D05CC341730F0F00C0FB0",
            INIT_RAM_26 => X"58A8990780D0A28AAABAEB057F44759B651054E090918885A69988304128C7D0",
            INIT_RAM_27 => X"849425411250A509B60C23A1D6CE8BBBBBB2A5A081039510825E6A49B2C612C0",
            INIT_RAM_28 => X"C4218C9F07B26C5128088424DB366822528884C4F257B15C813DCC4400882008",
            INIT_RAM_29 => X"8110050042A5A100AB2B282B8070743A4089FFFFF80A09C0012580E209D84820",
            INIT_RAM_2A => X"700686201F6926423EDC9480A506702617F4F4EDA4FAA449480A8056B4B23803",
            INIT_RAM_2B => X"24C3404309604B10854D05B902B2821021656808C29728050CB834D826C848C0",
            INIT_RAM_2C => X"46885301420A9939A842A6528463206B98D1A30909B0A861D012C21812CCAA14",
            INIT_RAM_2D => X"36A5816061BDD85296258186F72C3D1FE84FD4DCCFC2D1CD42994A918C85AE63",
            INIT_RAM_2E => X"48C442F0E1899FEE0016108C7FC5D020384135340815C4E92188823482AD9093",
            INIT_RAM_2F => X"3864735C89C9AA48FECF71211A303C3E3C343830C31FAD93A8C786BA3FD2F048",
            INIT_RAM_30 => X"21DBABB0908B584997B1989C936E98286828C1E84D50E58732B7905ACC2A468C",
            INIT_RAM_31 => X"656131A8B8576D8986CA046680C576C3DDD322EE0983DA1F0A8D1D681C80046A",
            INIT_RAM_32 => X"83C7852910A49C90421290C9138F1C551698E1C64981846824212077319A6069",
            INIT_RAM_33 => X"2002500385A0C78100110001243E8000EA46882236E47523400F0F65B48F0B93",
            INIT_RAM_34 => X"310731134AA556804442800C628A08201C40019F644800120225200441800628",
            INIT_RAM_35 => X"EA3F940E368260F809EA7FE24429A7FE28031E1048F08879C42049C090239848",
            INIT_RAM_36 => X"DB22117910FCCE77F557FFFFDD57F5757D7F5FFFD7F757FD5F5FF5F5FF400068",
            INIT_RAM_37 => X"093030E5EF7E2A0B0804DAC13B776198154409C6A33413E9230434AB4F355137",
            INIT_RAM_38 => X"021414662067C1AAAAAAA14021C60A1402142CB45EB44D4340240C8297248A98",
            INIT_RAM_39 => X"6969084198A0A12929C92928492949F90861802180F8719998092863FC9001B8",
            INIT_RAM_3A => X"3E0019F861F979E02061C101F92849484908706100F101F82108292909092849",
            INIT_RAM_3B => X"0BC01999F861728041E1810121501090911011E1F8E201E82290295121112150",
            INIT_RAM_3C => X"8C5CE06060639FB8C7CE5606063CDB8D7EE56060620538D7EE060600118D7EC0",
            INIT_RAM_3D => X"00000000006838C30C2006060041818181800060656063DFB881460656063DFB",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"4680000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"980CC6C1820883020862069D388E28E2098F29C4C67030600B00000201E800D3",
            INIT_RAM_01 => X"A13A220BB0610506080A4FA33EF8B88D0ABB8ECE11806860C00297DAFD3DF180",
            INIT_RAM_02 => X"4301D7C9D751820120A71893AA8C04423F5389E3B822E876A7FFFC0514AD0D6A",
            INIT_RAM_03 => X"6130181FFFE8C1247864D01B4E8A31461070CE5DCCA6110081FFE18065C10090",
            INIT_RAM_04 => X"6510980C0FFF04012E180C0A180EB6E4693AA8864D019068A714E1070CE5DCCA",
            INIT_RAM_05 => X"0B4A32852BFBEEDBB544406051A60102980C1820412280CA34538A70818672EE",
            INIT_RAM_06 => X"04880CC50AE38DFE902169059D1DC5FFC379E1B0F0484A62057BB288B820C110",
            INIT_RAM_07 => X"2C45227C1222DFBB9FFD95F72009297B9006ADA764086EF3A823F0E44935047E",
            INIT_RAM_08 => X"3F0244060202052AE3ADFE90214EBDEE93B3A3B8BFE82FA658065FFFE3FFD93F",
            INIT_RAM_09 => X"88B7EEE7FBE412B5411FFE84EC82492B20558301D3B2043779D411F872249A82",
            INIT_RAM_0A => X"321039EFF841C2146443FC860EB037E8B15930DF8017FFF8FFF6CFCB13489F04",
            INIT_RAM_0B => X"FC3FFF03FFE0AAAAAB94D1614A91900005E68F9BFE13C248FEA13D425F822012",
            INIT_RAM_0C => X"03FE8FB0627F0FFB89FDC0FF7EFE0807FD1F0313F844FFFFBC1FF7EFE1FFFFFF",
            INIT_RAM_0D => X"F1FC7FFF1F70FFE7F7CFFFE3EE1FFDFDFBEFEFA3EFD9FF8FF1FDBEF0C99FFFB8",
            INIT_RAM_0E => X"0956F1EC6318C6318C6318C6318FEFFDCFE7F7FB01C7FE73F7A3FE667EF0F9FF",
            INIT_RAM_0F => X"1E27E89251C28866ED9F750566B12CE506FBBB15078255812AC19560CABC12AC",
            INIT_RAM_10 => X"40686DDE01EC7C3C6005FA6B5A35D77CFF9326C9C4718BF491280C4337685116",
            INIT_RAM_11 => X"0745D400E8A85165C0AAF91F9324AAAE03F2BE9615F7F2A14C9287D5D644FD09",
            INIT_RAM_12 => X"0C8B0D56D230D871A2B105823D0F4B25208918380881C7EF92B111510888A89A",
            INIT_RAM_13 => X"1C130E03C149491482C8A86F1050C1608EABDDEAC176ECC3B0AC857211C76524",
            INIT_RAM_14 => X"4613C6B0AF88C192148C38F870ABEF9FAAA1832104A1AB4FFFFD1F21F20DA824",
            INIT_RAM_15 => X"FDFFFE07FE602200C75DB94E76B47168B9800C20692987806A77BA4CAAFFEA82",
            INIT_RAM_16 => X"38728C8993B568CE993362E5CA156EBAD7DFF89F1FFFFFE1EFF73FFC3FFDF41B",
            INIT_RAM_17 => X"F997DB3038DFBC0F441050154005500157FE3C7DEFA7EB446BFFE9E7D3F3E09C",
            INIT_RAM_18 => X"E92081171D156AB552A954AA401306DB090520781E0A9688348BDD7DC732E1DB",
            INIT_RAM_19 => X"730AD39FE617A60A2041966F80954217FD0DE9E9DC4A7605121B02D09140844B",
            INIT_RAM_1A => X"B6C5B6DB6D86DB6DB63FFFFFFCFFFE2282FFFA3BFFDE3BD20A262190E1C36C90",
            INIT_RAM_1B => X"FFC0F4F3FFF4FBD3FF4A7FFF4FD1F800000000003FFEFD861C18707FFFC2DB6D",
            INIT_RAM_1C => X"C3A1D0E8741A0F2244D558360096216283FFBBE3FF9F0460EFFFFDFFFFFC045F",
            INIT_RAM_1D => X"1FDE8FA1F60E8BD25A520401879A405E2C0448D97D7FD1B6EBD2C261D06C8908",
            INIT_RAM_1E => X"B5F8E46464095CB60104601B121588060E6019C1D6FD57BBB83DFBEEC1E04087",
            INIT_RAM_1F => X"44135047E04881CCEDBF6CFBB6F981D9D3DDBB6789EFDF7EFFF6FEFEFDEDF9EF",
            INIT_RAM_20 => X"F71FFD0FFD1085FF63885E15E08560AD24E67E437F6EC7C50B9106EF3A823F0E",
            INIT_RAM_21 => X"EDE67F35A2AB352A540AC7D66422E0AFA373DBE4707AC1FA2C7748E4029933FF",
            INIT_RAM_22 => X"D123A247460CF0FBEDFDBFB7F6FADF5BEB7D6F7DF6FADF5BEB7F6FEDFDBFB7BD",
            INIT_RAM_23 => X"D35DFF7FF9FFFF6C6AF1086C70404D181820F00B06715D04622C384C1C1E8991",
            INIT_RAM_24 => X"80C3017E815C6B1057E832C7DDF20AE432C60EA230AC53E0AE9142F1F2A8F8BF",
            INIT_RAM_25 => X"F87FE1EE08ECACD8EB577642077B696429308D1A2F9FD7FC7F5FF1F1F1FF807B",
            INIT_RAM_26 => X"FB2981FAFAFF5965144105F8879E5A0857EAAF0760014F10DD41F77107FB8037",
            INIT_RAM_27 => X"1D9D6711846046039E620B65A02D907E5A18032186C42B70C70540E907C80502",
            INIT_RAM_28 => X"08518FA038503CCA6A652526A08FC194D7E535B215C88A78627A028408C232CE",
            INIT_RAM_29 => X"F75DDDDDD7DDF75F7BFBFA1FF979FF05035E08282092EB5240FF43EFE1E32571",
            INIT_RAM_2A => X"09FDFDFF8087FDFF01005B27EC255142B019435A84B36085F807FFFFF8EE97BB",
            INIT_RAM_2B => X"34D7035E2AC2160504D81F765F958AB140AFC8FCE4AD582885F742405F94C406",
            INIT_RAM_2C => X"A59FC20E619743413C7DCD7E4CD612F889E96579F421442B80D78AF085856828",
            INIT_RAM_2D => X"7165594448F9F41595651123E7CCADAE300023B69DD53709E335F9B3584BE227",
            INIT_RAM_2E => X"00A68878F1F41FFF71E08388E03292A38D9F0CA47DB3B355B514361B25E05B90",
            INIT_RAM_2F => X"FDEBFB7D81E1D483D58911631E3D6B256F276F2CDFBDBD270C628A16755D02B0",
            INIT_RAM_30 => X"CFFBCAF0ED8E9EACE831C86EFA8F82445438F0047D17CB07963D7479C405458A",
            INIT_RAM_31 => X"C2C314403C3D7B9BA7EA4458538154D291F04788F247A10B17895CC60F8FFFFF",
            INIT_RAM_32 => X"87E9BFBC8574BF4A22195EAD5625A0181715F080730B0A993DEF652D2014CAC6",
            INIT_RAM_33 => X"CC5FFF90E37D002FFDFEFFFF7E0FFFE3EFFFDEBFFFFDF7FFEFFF07FB5F404252",
            INIT_RAM_34 => X"11FAF7AFFD7AF77BE998F98C628A3FFFF8037F00FDFFEBFFF9FFFF87F60758C7",
            INIT_RAM_35 => X"F638FDFFBF7FFFFFF017B81FFFFBC0026B30ABFF855FFC07F87D7F3BF87FFFFC",
            INIT_RAM_36 => X"FDFFFFFE01F9FFDD5557FFFD5FFD557FD57FF55FFD57FD555FF555FF554803F0",
            INIT_RAM_37 => X"C7FFDFB7FFFDFFDF47FF83FFFFFFBFEEFA7FF5FF011F03FDBF7FBFFFFF1FFFFD",
            INIT_RAM_38 => X"020154667BBF8FFFFFFFFFFFF7F7DFFFFF7FFFF87FE99EFEFDFF7FFFDEFFF7FF",
            INIT_RAM_39 => X"08080040F1A00129298939285909C9F988C000210020E108F001F8D129F80000",
            INIT_RAM_3A => X"1E00310831F9E9E070C0E101F928490849083831006101082198292909992859",
            INIT_RAM_3B => X"0B8009080001F280E100C101F950109091101010F84201E82293F95121112150",
            INIT_RAM_3C => X"0E79C0604043BFF0E7DC5604043FFF0F7FC52040439A70F7FC040439A7077EC0",
            INIT_RAM_3D => X"000000000042B082082204043DA90101010F7A40650043FFF077AC0654043FFF",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"402A04C5405401150110024588C60C60450F0543318DCF9FFC0101010017F7B1",
            INIT_RAM_01 => X"40C9512610082A005404AFA29E510044411784950AC2B39F3FFD5FFA5D35F024",
            INIT_RAM_02 => X"9A829A254E0AB50AC1112B58EEC422011F1A8D61C8A148D0C000020144E224B0",
            INIT_RAM_03 => X"50A854239CE55A9FF1161810627B11621151FC8520910A854039AC4313988460",
            INIT_RAM_04 => X"04A8542A01CD6A1A9CC42214C414D11224AEFF95698122A7B11621111FC85209",
            INIT_RAM_05 => X"0E5FFB057A2D286A1882A11008910884442A01108AB4C09353D88B10888FE429",
            INIT_RAM_06 => X"43FB80C8BC2F35FED802F00E859B8EF60AECC428C214460603CA1A0799100880",
            INIT_RAM_07 => X"0E01B9569B91DB6D01FAB46192601B70C937CBC38025023D1C6EB2DFED638DD6",
            INIT_RAM_08 => X"EB01FDC01504C89C2F15FED802FE1C9702D0B373DED15DC200030FFBDDF7F81A",
            INIT_RAM_09 => X"E476DB5077E80A18E375FD14264285A990794A82E1C012811E8E37586FF6B1C6",
            INIT_RAM_0A => X"1E20509002C840030A026A110A464A40EC1EE2BCA043FEF77DFE0683806E45A6",
            INIT_RAM_0B => X"DFFFFFE014008200830931A8E1C297FFE6E5190D29192311295192A31081108C",
            INIT_RAM_0C => X"00DF77C19D8FC03C763E0F00BF7F8C01BEEF8CEC7E3B1F7FC0E00BF7F9FDB7FD",
            INIT_RAM_0D => X"EEFE1FBEEFBC001BF803F7DDF780FEFEFC03F7DDF7E8FF77DBFEDF08306003DE",
            INIT_RAM_0E => X"44000E0318C6318C6318C6318C60701E77F00B7CFE27F18CFBD3F9999F7C06DF",
            INIT_RAM_0F => X"06A03FCA107BF072065A318064208E29CCD731DF8795000A80044002200C8800",
            INIT_RAM_10 => X"4F70640E2FB9B5F4DD82A8DA5C65D74872B9738D46B0F01E7D09EF8390351206",
            INIT_RAM_11 => X"414C450C298A76BAC09E9032B9702D5E009AFF4249A3189468DE54499A9404D8",
            INIT_RAM_12 => X"1508117B4B58501A9EF54CCC86FF45ADB457067A1943DCA4D262AAA9F15554E4",
            INIT_RAM_13 => X"688D7A1FCC60EF0C018095A4622088C053234DA0CAB26D40803C01E1188266D8",
            INIT_RAM_14 => X"1E1AC3007D08C294038C087813F9659FF9E4814082610543FC34AFD2FD0A00B2",
            INIT_RAM_15 => X"FEBFCF80FF1FDDFF2C9F9B6EA4B8A57150201899CC8F3CB7A5908B6B99C3EE59",
            INIT_RAM_16 => X"DBA54B0E9C2950B2E9D2852A542A104130C3FEC08FE2FEF8000B8FFF03FE7BE3",
            INIT_RAM_17 => X"FB15D824B0CFBC0F461500155550000151FDC38C17DBF439000FF01BF80DF969",
            INIT_RAM_18 => X"D5B74C212F273B9FCFE773B9ED6E16013100B7F9FE2E4CD9140FD97D4210E2A0",
            INIT_RAM_19 => X"7633578AA56DB5212B2722E50219D93154A725654C2426BF19735954C1E19394",
            INIT_RAM_1A => X"496649249249249249000000007EFF1D7C0001FC3FE1FF9619D99370A142CDA2",
            INIT_RAM_1B => X"7FE0FC13E1FCFDF07FC61FDFC5F0FD7C1F003E0F9EDF1E082220883F7FC36492",
            INIT_RAM_1C => X"4A8542A150A855428340088CC2C10102483BCC1003C0FB9F03FDFC7DEF7F02A3",
            INIT_RAM_1D => X"87EF43DE090F744DCDCE5B6447BB0B3428124098D8DBD937FFD281C442250A04",
            INIT_RAM_1E => X"CCA9B0303064F7DAB0622208100D0B04132E0C82D23F30889800FDF7381FBF78",
            INIT_RAM_1F => X"FED638DD643FB989B4DD3C26D370C0302166EDE64470078001FB7F001EF6FE03",
            INIT_RAM_20 => X"7B801E01BEE7829A84506216208E204558383281C9B3725A07E25133D1C6EB2D",
            INIT_RAM_21 => X"1203BFE5C54172244818CD22C16620021E4D7350A829189033AEA11C10460C00",
            INIT_RAM_22 => X"A0E141C281038000120640C8190720E41C839000090720E41C8390720E41C802",
            INIT_RAM_23 => X"507F862FFC71C9241A8CE78CD831B2E486196D5D3CF4625411820A121E0D0C70",
            INIT_RAM_24 => X"7F2E02FF61AC3012AF52F795C85E55E810020E1FBA0EAFF15EDAA5F359F9E81F",
            INIT_RAM_25 => X"FE7FFBEDA05B5B68020E06EA5A1656371FAA97101000280200A00808087FE000",
            INIT_RAM_26 => X"7870647EF51FCF3CF3DF7DFF87EFD284CD01418ACC2C62808E240B88E03C60E7",
            INIT_RAM_27 => X"FC73BDE73BDE3DE7BF358311980C4D979A68FBA18763BC8E3204032A92518020",
            INIT_RAM_28 => X"380DAC7E57F07C859CB2CF2471BAC6CB7AB2DED9D37D85C8313F417DC7BDEF39",
            INIT_RAM_29 => X"381EE1EE07E1F81F800000EFBC3C3FFF238FF775D54A532EB9FFBC10FD459630",
            INIT_RAM_2A => X"06FE1C7FC07B7C7F80F034C8B2CE72211A90505C32FAA4430CBBEF7FBCF02BC0",
            INIT_RAM_2B => X"069A026A2D422A1A85658191225881122115642B4AD5A854023989240C8C0C09",
            INIT_RAM_2C => X"E30A2F15002B24B7A857FEFB17F08C6CCBB8C1A95262A01500988B1088822A54",
            INIT_RAM_2D => X"F3318C6A9134D3044611AA44D314BD162E601DFCDD82DCBD43FBEC5FC031B22E",
            INIT_RAM_2E => X"1630404081124007B81F78CE601CDB0018C192740898DA4A21889E10C8B230EC",
            INIT_RAM_2F => X"2840D61A7743AB62568C50230A28F4F0F0F0F0F38D1E6501ABB2A601A80A4466",
            INIT_RAM_30 => X"2B4AA092C966249816F088430C1A65D2627880126D0243820211047BC418C080",
            INIT_RAM_31 => X"1010E0B7A81C3904489C04292D101E93C30CBF3A098EE4932CDC17F40860F7FC",
            INIT_RAM_32 => X"F2E104E602BBDC25920024B623AE5BD6CA91A1C68840448080002146F1A21410",
            INIT_RAM_33 => X"E3837F281DBEF043EEF6EFBFBF87BFD0F37F8143BEFC79BFC7BFC87DA7A0A375",
            INIT_RAM_34 => X"287E3BE3CCBE191C7AA8024E73CF0EFDFBF0BFC0247FF01FFC7DFCE009E0063B",
            INIT_RAM_35 => X"79981EE0406FF7FEFC0BD803FDFDF0018448D781E6BC1F01F7028CDCFE0001FF",
            INIT_RAM_36 => X"1FFFFFFFFFE7FFEAAAA800000AAAAA80002AAAA00002AAAAA00000AAAAA7F1FC",
            INIT_RAM_37 => X"FFFFFFC80002FFEFB8077FFF7FF84FFF7DFEFE3FFEFFFFFEFFBFFFFFFFFFDDFE",
            INIT_RAM_38 => X"02555419FFFFF7E00001EFDBFFFFFEFDBFFF841783F66FFFDFFFFFFFFF3DFFFF",
            INIT_RAM_39 => X"F818004061000139F809F1B87199D910F18000200020A0006000D1A939F83800",
            INIT_RAM_3A => X"0E0021081801C839D9F879F809B9F9F9F9F9F9F9F9F98109F8F1F9F9F8F1F9F1",
            INIT_RAM_3B => X"0B0010000001D2F1B1F071F0F971E0F3F1F1E1F001FB0001FAF3F1F1E1F1F9D0",
            INIT_RAM_3C => X"0A3580200000EDE0A3585200000EDC0B37852000008D403378000008500337A0",
            INIT_RAM_3D => X"000000000040308249220000241C000000010600250000EDE091700250000EDE",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"FF80000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"406A048548560315215802D4A8544564D5050C40000000000C010103000002D1",
            INIT_RAM_01 => X"E089110630006B00D4042EA00AE010550112808418C238000004555A5515706C",
            INIT_RAM_02 => X"8A870C455A0A951A8035738AAA546A0355488465D02000724000028050601480",
            INIT_RAM_03 => X"11A8D42308CD5AB7515688126A2B506A0110EC892435188C4231C44316888C40",
            INIT_RAM_04 => X"2188D46A118E2A1ABC546A1054386522A48AAE9160800222B10620110EC89243",
            INIT_RAM_05 => X"0E53AB803A2B287A1C8623501AB51A80D462035008B040831158831008876449",
            INIT_RAM_06 => X"115340C8B44539FE4882E81A888A9A0A18ACEC08D684431203D21A029B101880",
            INIT_RAM_07 => X"060099528991C96542F9B09232405B091924838300A504510A2B884AAD614571",
            INIT_RAM_08 => X"B8A0A9A0350448B44739FE4802EE9D8E8251137141C31DA2081300000000181E",
            INIT_RAM_09 => X"6476D940AFF01218515C7CB442C014A0B0105882C1805282288515C56556B0A2",
            INIT_RAM_0A => X"0A0010900098A0214A02C93502560A402810863D2100000000060783802644A2",
            INIT_RAM_0B => X"0001400014000000010935E9E3C752AAA7619A4F49592B01495192A301131188",
            INIT_RAM_0C => X"00000004000020000000000000004A0000002000010000000000000004000000",
            INIT_RAM_0D => X"0000000000020000000000000040000000000000000C00000000000000000001",
            INIT_RAM_0E => X"4402000000000000000000000000000000000000001000000008000000020000",
            INIT_RAM_0F => X"04801542008B58520240338040608E41CC85205A8591008880444022201C8804",
            INIT_RAM_10 => X"094844062D09A1A05987005A5E655752749933844232E00A2900AAC290151604",
            INIT_RAM_11 => X"424C8508498A508EC0BEA43499322FF6008ADA021C03380048DF14C33C100018",
            INIT_RAM_12 => X"0408115FD950401ABBB54C5D93D746AC945F043A0941DD04D042AAA8E155546E",
            INIT_RAM_13 => X"718D6A15C420EF0A03D080A426B09A8055224CA098B26542802C0173088A46DC",
            INIT_RAM_14 => X"0E0ACB203C08C090038C087813F9C716F8E4814086E10F0B780DA01A01820016",
            INIT_RAM_15 => X"000020DE000000011CD49B68A4BCA579D0A019BBC5871D33A5C21123B343E6CB",
            INIT_RAM_16 => X"E3E78FEFDF3F78FEFDFBD7AF1E3F7EEBF7D8018C401800042000000080020004",
            INIT_RAM_17 => X"FB111014306B940944000015555555540000004C000002046A000000120005F9",
            INIT_RAM_18 => X"94944402050A150A84422110880E0601010992A8AE66DC93140D4D3DC2304084",
            INIT_RAM_19 => X"6233C7A0052D9503692716A2001DC930008724644C04249E097249D001A1B794",
            INIT_RAM_1A => X"001800000030000000C00000030000800000000000000396199990702040C982",
            INIT_RAM_1B => X"000F07FC1007041F007FC0007C1E02FFE00001FF80000171C1C70780007C0000",
            INIT_RAM_1C => X"5A8D46A351A8D742831559ACC6450102D800201800000000000003000000FE00",
            INIT_RAM_1D => X"4000A00002B00045CDCECB25429B19702836409078794126E942836C46250A0C",
            INIT_RAM_1E => X"3C01E060606DE7DEB0666248101D0B86032E0CC05683FFFFFFFC000004000000",
            INIT_RAM_1F => X"AAD6145710153489906D1CA641B0423235230626450090040000000000000208",
            INIT_RAM_20 => X"00000000000482920D506A06A00EA0D420103481D0C1929007DA504510A2B88C",
            INIT_RAM_21 => X"00000065E540502040108120804E40005B0C7649882958900AA4011430400000",
            INIT_RAM_22 => X"A06140C28321A000000C0180300600C018030000000200400801002004008000",
            INIT_RAM_23 => X"C2FF01600100096DFAAC42C8C81126ACA208441C3674765530860A161E0D0C30",
            INIT_RAM_24 => X"001B00DF60ACB210AD527795409E15A010420E1EA208AAE15A4A21B218F9B81F",
            INIT_RAM_25 => X"010006ADA05B5B78020424CC5A1316B717A31610000800052000149494001FF8",
            INIT_RAM_26 => X"2A506D070C007FFFFFFFFE03F820D28DDC011198CC642080AF6C1805D400D7F0",
            INIT_RAM_27 => X"5CD694AD694A14A3AB14C6130918453D9278CA2107336CCA1604006802918221",
            INIT_RAM_28 => X"380D0C7E57E0148CB4B65B0028AE10D928364A5BD33D8CD21937433546B4A529",
            INIT_RAM_29 => X"0000000000000000000000000000007F23AFE280AC0012249000000005C7B232",
            INIT_RAM_2A => X"F0004200BFFB02017FF874CAB25F66A35A90505E36DC24474C80000000000000",
            INIT_RAM_2B => X"020A026A0D402A0A802585222A4A8156A0312C098C4488C4063DDB640D86240E",
            INIT_RAM_2C => X"33082735002B6C93A047EA69189205640988C08916E6203180188310088620C4",
            INIT_RAM_2D => X"FB31CC6A98D0D304C731AA6341381D53FD5FFCFCD480DC9D03A9A4E24A119126",
            INIT_RAM_2E => X"32104050A156C000000005AD3FFDC9411AC482F42A894A499C8C0C54C8B074ED",
            INIT_RAM_2F => X"2840961A7302AB62978C50A30A2070F070F070FB8D1A6901ABE084418A224C66",
            INIT_RAM_30 => X"3F52AAA0C966240C567088034D386DD67658803635028382021114394411C080",
            INIT_RAM_31 => X"3838E833201D3B42CAB4040B6F300E93C70DB7186004AD920C9013B00A600002",
            INIT_RAM_32 => X"D08344E706BB4D6DB2002C9BB00AD996589101C7A8E0E48C84219852F1EA3838",
            INIT_RAM_33 => X"085800B740000FE0020100008070002A00004000000500002001A000005FE361",
            INIT_RAM_34 => X"B50780384F83C1C00FFACBAD6BAEA00007E8803FE50018C00700021300177080",
            INIT_RAM_35 => X"004F00000180000003F80FE000040FFC6F770044180240FC0000000001000000",
            INIT_RAM_36 => X"010408011112100AAAAAAAAAA0000000002AAAAAAAA80000000000AAAAA00802",
            INIT_RAM_37 => X"24101020210A0000040482020114000800400520491042012200200220908021",
            INIT_RAM_38 => X"0200004442204815555500000404100000404104820888808100402210800408",
            INIT_RAM_39 => X"F010000000000010D008E0B86091910061000000000000000000011010901800",
            INIT_RAM_3A => X"060000000801881999F838F80891F8F1F8F1F9F9F9F88001F861F9F9F861F9E0",
            INIT_RAM_3B => X"0A0000000001927110F030F00021F063F0E1F1E001F90001F86000E0C0E1F880",
            INIT_RAM_3C => X"0F638000000178E0F6385000001F8E077F85000001D8E073FA0000358E073F80",
            INIT_RAM_3D => X"000000000055528A28A80000154A008000075380050000E8E0F6380050000E0E",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

end Behavioral; --Gowin_pROM
